/* modified netlist. Source: module Asconp in file ./test/Asconp.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

// `include "General/Gates.v"

module Asconp_HPC2_ClockGating_d1 (state_in_s0, rcon, clk, state_in_s1, Fresh, /*rst,*/ state_out_s0, state_out_s1/*, Synch*/);
    input [319:0] state_in_s0 ;
    input [3:0] rcon ;
    input clk ;
    input [319:0] state_in_s1 ;
    //input rst ;
    input [319:0] Fresh ;
    output [319:0] state_out_s0 ;
    output [319:0] state_out_s1 ;
    //output Synch ;
    wire n3230 ;
    wire n3231 ;
    wire n3232 ;
    wire n3233 ;
    wire n3234 ;
    wire n3235 ;
    wire n3236 ;
    wire n3237 ;
    wire n3238 ;
    wire n3239 ;
    wire n3240 ;
    wire n3241 ;
    wire n3242 ;
    wire n3243 ;
    wire n3244 ;
    wire n3245 ;
    wire n3246 ;
    wire n3247 ;
    wire n3248 ;
    wire n3249 ;
    wire n3250 ;
    wire n3251 ;
    wire n3252 ;
    wire n3253 ;
    wire n3254 ;
    wire n3255 ;
    wire n3256 ;
    wire n3257 ;
    wire n3258 ;
    wire n3259 ;
    wire n3260 ;
    wire n3261 ;
    wire n3262 ;
    wire n3263 ;
    wire n3264 ;
    wire n3265 ;
    wire n3266 ;
    wire n3267 ;
    wire n3268 ;
    wire n3269 ;
    wire n3270 ;
    wire n3271 ;
    wire n3272 ;
    wire n3273 ;
    wire n3274 ;
    wire n3275 ;
    wire n3276 ;
    wire n3277 ;
    wire n3278 ;
    wire n3279 ;
    wire n3280 ;
    wire n3281 ;
    wire n3282 ;
    wire n3283 ;
    wire n3284 ;
    wire n3285 ;
    wire n3286 ;
    wire n3287 ;
    wire n3288 ;
    wire n3289 ;
    wire n3290 ;
    wire n3291 ;
    wire n3292 ;
    wire n3293 ;
    wire n3294 ;
    wire n3295 ;
    wire n3296 ;
    wire n3297 ;
    wire n3298 ;
    wire n3299 ;
    wire n3300 ;
    wire n3301 ;
    wire n3302 ;
    wire n3303 ;
    wire n3304 ;
    wire n3305 ;
    wire n3306 ;
    wire n3307 ;
    wire n3308 ;
    wire n3309 ;
    wire n3310 ;
    wire n3311 ;
    wire n3312 ;
    wire n3313 ;
    wire n3314 ;
    wire n3315 ;
    wire n3316 ;
    wire n3317 ;
    wire n3318 ;
    wire n3319 ;
    wire n3320 ;
    wire n3321 ;
    wire n3322 ;
    wire n3323 ;
    wire n3324 ;
    wire n3325 ;
    wire n3326 ;
    wire n3327 ;
    wire n3328 ;
    wire n3329 ;
    wire n3330 ;
    wire n3331 ;
    wire n3332 ;
    wire n3333 ;
    wire n3334 ;
    wire n3335 ;
    wire n3336 ;
    wire n3337 ;
    wire n3338 ;
    wire n3339 ;
    wire n3340 ;
    wire n3341 ;
    wire n3342 ;
    wire n3343 ;
    wire n3344 ;
    wire n3345 ;
    wire n3346 ;
    wire n3347 ;
    wire n3348 ;
    wire n3349 ;
    wire n3350 ;
    wire n3351 ;
    wire n3352 ;
    wire n3353 ;
    wire n3354 ;
    wire n3355 ;
    wire n3356 ;
    wire n3357 ;
    wire n3358 ;
    wire n3359 ;
    wire n3360 ;
    wire n3361 ;
    wire n3362 ;
    wire n3363 ;
    wire n3364 ;
    wire n3365 ;
    wire n3366 ;
    wire n3367 ;
    wire n3368 ;
    wire n3369 ;
    wire n3370 ;
    wire n3371 ;
    wire n3372 ;
    wire n3373 ;
    wire n3374 ;
    wire n3375 ;
    wire n3376 ;
    wire n3377 ;
    wire n3378 ;
    wire n3379 ;
    wire n3380 ;
    wire n3381 ;
    wire n3382 ;
    wire n3383 ;
    wire n3384 ;
    wire n3385 ;
    wire n3386 ;
    wire n3387 ;
    wire n3388 ;
    wire n3389 ;
    wire n3390 ;
    wire n3391 ;
    wire n3392 ;
    wire n3393 ;
    wire n3394 ;
    wire n3395 ;
    wire n3396 ;
    wire n3397 ;
    wire n3398 ;
    wire n3399 ;
    wire n3400 ;
    wire n3401 ;
    wire n3402 ;
    wire n3403 ;
    wire n3404 ;
    wire n3405 ;
    wire n3406 ;
    wire n3407 ;
    wire n3408 ;
    wire n3409 ;
    wire n3410 ;
    wire n3411 ;
    wire n3412 ;
    wire n3413 ;
    wire n3414 ;
    wire n3415 ;
    wire n3416 ;
    wire n3417 ;
    wire n3418 ;
    wire n3419 ;
    wire n3420 ;
    wire n3421 ;
    wire n3422 ;
    wire n3423 ;
    wire n3424 ;
    wire n3425 ;
    wire n3426 ;
    wire n3427 ;
    wire n3428 ;
    wire n3429 ;
    wire n3430 ;
    wire n3431 ;
    wire n3432 ;
    wire n3433 ;
    wire n3434 ;
    wire n3435 ;
    wire n3436 ;
    wire n3437 ;
    wire n3438 ;
    wire n3439 ;
    wire n3440 ;
    wire n3441 ;
    wire n3442 ;
    wire n3443 ;
    wire n3444 ;
    wire n3445 ;
    wire n3446 ;
    wire n3447 ;
    wire n3448 ;
    wire n3449 ;
    wire n3450 ;
    wire n3451 ;
    wire n3452 ;
    wire n3453 ;
    wire n3454 ;
    wire n3455 ;
    wire n3456 ;
    wire n3457 ;
    wire n3458 ;
    wire n3459 ;
    wire n3460 ;
    wire n3461 ;
    wire n3462 ;
    wire n3463 ;
    wire n3464 ;
    wire n3465 ;
    wire n3466 ;
    wire n3467 ;
    wire n3468 ;
    wire n3469 ;
    wire n3470 ;
    wire n3471 ;
    wire n3472 ;
    wire n3473 ;
    wire n3474 ;
    wire n3475 ;
    wire n3476 ;
    wire n3477 ;
    wire n3478 ;
    wire n3479 ;
    wire n3480 ;
    wire n3481 ;
    wire n3482 ;
    wire n3483 ;
    wire n3484 ;
    wire n3485 ;
    wire n3486 ;
    wire n3487 ;
    wire n3488 ;
    wire n3489 ;
    wire n3490 ;
    wire n3491 ;
    wire n3492 ;
    wire n3493 ;
    wire n3494 ;
    wire n3495 ;
    wire n3496 ;
    wire n3497 ;
    wire n3498 ;
    wire n3499 ;
    wire n3500 ;
    wire n3501 ;
    wire n3502 ;
    wire n3503 ;
    wire n3504 ;
    wire n3505 ;
    wire n3506 ;
    wire n3507 ;
    wire n3508 ;
    wire n3509 ;
    wire n3510 ;
    wire n3511 ;
    wire n3512 ;
    wire n3513 ;
    wire n3514 ;
    wire n3515 ;
    wire n3516 ;
    wire n3517 ;
    wire n3518 ;
    wire n3519 ;
    wire n3520 ;
    wire n3521 ;
    wire n3522 ;
    wire n3523 ;
    wire n3524 ;
    wire n3525 ;
    wire n3526 ;
    wire n3527 ;
    wire n3528 ;
    wire n3529 ;
    wire n3530 ;
    wire n3531 ;
    wire n3532 ;
    wire n3533 ;
    wire n3534 ;
    wire n3535 ;
    wire n3536 ;
    wire n3537 ;
    wire n3538 ;
    wire n3539 ;
    wire n3540 ;
    wire n3541 ;
    wire n3542 ;
    wire n3543 ;
    wire n3544 ;
    wire n3545 ;
    wire n3546 ;
    wire n3547 ;
    wire n3548 ;
    wire n3549 ;
    wire n3550 ;
    wire n3551 ;
    wire n3552 ;
    wire n3553 ;
    wire n3554 ;
    wire n3555 ;
    wire n3556 ;
    wire n3557 ;
    wire n3558 ;
    wire n3559 ;
    wire n3560 ;
    wire n3561 ;
    wire n3562 ;
    wire n3563 ;
    wire n3564 ;
    wire n3565 ;
    wire n3566 ;
    wire n3567 ;
    wire n3568 ;
    wire n3569 ;
    wire n3570 ;
    wire n3571 ;
    wire n3572 ;
    wire n3573 ;
    wire n3574 ;
    wire n3575 ;
    wire n3576 ;
    wire n3577 ;
    wire n3578 ;
    wire n3579 ;
    wire n3580 ;
    wire n3581 ;
    wire n3582 ;
    wire n3583 ;
    wire n3584 ;
    wire n3585 ;
    wire n3586 ;
    wire n3587 ;
    wire n3588 ;
    wire n3589 ;
    wire n3590 ;
    wire n3591 ;
    wire n3592 ;
    wire n3593 ;
    wire n3594 ;
    wire n3595 ;
    wire n3596 ;
    wire n3597 ;
    wire n3598 ;
    wire n3599 ;
    wire n3600 ;
    wire n3601 ;
    wire n3602 ;
    wire n3603 ;
    wire n3604 ;
    wire n3605 ;
    wire n3606 ;
    wire n3607 ;
    wire n3608 ;
    wire n3609 ;
    wire n3610 ;
    wire n3611 ;
    wire n3612 ;
    wire n3613 ;
    wire n3614 ;
    wire n3615 ;
    wire n3616 ;
    wire n3617 ;
    wire n3618 ;
    wire n3619 ;
    wire n3620 ;
    wire n3621 ;
    wire n3622 ;
    wire n3623 ;
    wire n3624 ;
    wire n3625 ;
    wire n3626 ;
    wire n3627 ;
    wire n3628 ;
    wire n3629 ;
    wire n3630 ;
    wire n3631 ;
    wire n3632 ;
    wire n3633 ;
    wire n3634 ;
    wire n3635 ;
    wire n3636 ;
    wire n3637 ;
    wire n3638 ;
    wire n3639 ;
    wire n3640 ;
    wire n3641 ;
    wire n3642 ;
    wire n3643 ;
    wire n3644 ;
    wire n3645 ;
    wire n3646 ;
    wire n3647 ;
    wire n3648 ;
    wire n3649 ;
    wire n3650 ;
    wire n3651 ;
    wire n3652 ;
    wire n3653 ;
    wire n3654 ;
    wire n3655 ;
    wire n3656 ;
    wire n3657 ;
    wire n3658 ;
    wire n3659 ;
    wire n3660 ;
    wire n3661 ;
    wire n3662 ;
    wire n3663 ;
    wire n3664 ;
    wire n3665 ;
    wire n3666 ;
    wire n3667 ;
    wire n3668 ;
    wire n3669 ;
    wire n3670 ;
    wire n3671 ;
    wire n3672 ;
    wire n3673 ;
    wire n3674 ;
    wire n3675 ;
    wire n3676 ;
    wire n3677 ;
    wire n3678 ;
    wire n3679 ;
    wire n3680 ;
    wire n3681 ;
    wire n3682 ;
    wire n3683 ;
    wire n3684 ;
    wire n3685 ;
    wire n3686 ;
    wire n3687 ;
    wire n3688 ;
    wire n3689 ;
    wire n3690 ;
    wire n3691 ;
    wire n3692 ;
    wire n3693 ;
    wire n3694 ;
    wire n3695 ;
    wire n3696 ;
    wire n3697 ;
    wire n3698 ;
    wire n3699 ;
    wire n3700 ;
    wire n3701 ;
    wire n3702 ;
    wire n3703 ;
    wire n3704 ;
    wire n3705 ;
    wire n3706 ;
    wire n3707 ;
    wire n3708 ;
    wire n3709 ;
    wire n3710 ;
    wire n3711 ;
    wire n3712 ;
    wire n3713 ;
    wire n3714 ;
    wire n3715 ;
    wire n3716 ;
    wire n3717 ;
    wire n3718 ;
    wire n3719 ;
    wire n3720 ;
    wire n3721 ;
    wire n3722 ;
    wire n3723 ;
    wire n3724 ;
    wire n3725 ;
    wire n3726 ;
    wire n3727 ;
    wire n3728 ;
    wire n3729 ;
    wire n3730 ;
    wire n3731 ;
    wire n3732 ;
    wire n3733 ;
    wire n3734 ;
    wire n3735 ;
    wire n3736 ;
    wire n3737 ;
    wire n3738 ;
    wire n3739 ;
    wire n3740 ;
    wire n3741 ;
    wire n3742 ;
    wire n3743 ;
    wire n3744 ;
    wire n3745 ;
    wire n3746 ;
    wire n3747 ;
    wire n3748 ;
    wire n3749 ;
    wire n3750 ;
    wire n3751 ;
    wire n3752 ;
    wire n3753 ;
    wire n3754 ;
    wire n3755 ;
    wire n3756 ;
    wire n3757 ;
    wire n3758 ;
    wire n3759 ;
    wire n3760 ;
    wire n3761 ;
    wire n3762 ;
    wire n3763 ;
    wire n3764 ;
    wire n3765 ;
    wire n3766 ;
    wire n3767 ;
    wire n3768 ;
    wire n3769 ;
    wire n3770 ;
    wire n3771 ;
    wire n3772 ;
    wire n3773 ;
    wire n3774 ;
    wire n3775 ;
    wire n3776 ;
    wire n3777 ;
    wire n3778 ;
    wire n3779 ;
    wire n3780 ;
    wire n3781 ;
    wire n3782 ;
    wire n3783 ;
    wire n3784 ;
    wire n3785 ;
    wire n3786 ;
    wire n3787 ;
    wire n3788 ;
    wire n3789 ;
    wire n3790 ;
    wire n3791 ;
    wire n3792 ;
    wire n3793 ;
    wire n3794 ;
    wire n3795 ;
    wire n3796 ;
    wire n3797 ;
    wire n3798 ;
    wire n3799 ;
    wire n3800 ;
    wire n3801 ;
    wire n3802 ;
    wire n3803 ;
    wire n3804 ;
    wire n3805 ;
    wire n3806 ;
    wire n3807 ;
    wire n3808 ;
    wire n3809 ;
    wire n3810 ;
    wire n3811 ;
    wire n3812 ;
    wire n3813 ;
    wire n3814 ;
    wire n3815 ;
    wire n3816 ;
    wire n3817 ;
    wire n3818 ;
    wire n3819 ;
    wire n3820 ;
    wire n3821 ;
    wire n3822 ;
    wire n3823 ;
    wire n3824 ;
    wire n3825 ;
    wire n3826 ;
    wire n3827 ;
    wire n3828 ;
    wire n3829 ;
    wire n3830 ;
    wire n3831 ;
    wire n3832 ;
    wire n3833 ;
    wire n3834 ;
    wire n3835 ;
    wire n3836 ;
    wire n3837 ;
    wire n3838 ;
    wire n3839 ;
    wire n3840 ;
    wire n3841 ;
    wire n3842 ;
    wire n3843 ;
    wire n3844 ;
    wire n3845 ;
    wire n3846 ;
    wire n3847 ;
    wire n3848 ;
    wire n3849 ;
    wire n3850 ;
    wire n3851 ;
    wire n3852 ;
    wire n3853 ;
    wire n3854 ;
    wire n3855 ;
    wire n3856 ;
    wire n3857 ;
    wire n3858 ;
    wire n3859 ;
    wire n3860 ;
    wire n3861 ;
    wire n3862 ;
    wire n3863 ;
    wire n3864 ;
    wire n3865 ;
    wire n3866 ;
    wire n3867 ;
    wire n3868 ;
    wire n3869 ;
    wire n3870 ;
    wire n3871 ;
    wire n3872 ;
    wire n3873 ;
    wire n3874 ;
    wire n3875 ;
    wire n3876 ;
    wire n3877 ;
    wire n3878 ;
    wire n3879 ;
    wire n3880 ;
    wire n3881 ;
    wire n3882 ;
    wire n3883 ;
    wire n3884 ;
    wire n3885 ;
    wire n3886 ;
    wire n3887 ;
    wire n3888 ;
    wire n3889 ;
    wire n3890 ;
    wire n3891 ;
    wire n3892 ;
    wire n3893 ;
    wire n3894 ;
    wire n3895 ;
    wire n3896 ;
    wire n3897 ;
    wire n3898 ;
    wire n3899 ;
    wire n3900 ;
    wire n3901 ;
    wire n3902 ;
    wire n3903 ;
    wire n3904 ;
    wire n3905 ;
    wire n3906 ;
    wire n3907 ;
    wire n3908 ;
    wire n3909 ;
    wire n3910 ;
    wire n3911 ;
    wire n3912 ;
    wire n3913 ;
    wire n3914 ;
    wire n3915 ;
    wire n3916 ;
    wire n3917 ;
    wire n3918 ;
    wire n3919 ;
    wire n3920 ;
    wire n3921 ;
    wire n3922 ;
    wire n3923 ;
    wire n3924 ;
    wire n3925 ;
    wire n3926 ;
    wire n3927 ;
    wire n3928 ;
    wire n3929 ;
    wire n3930 ;
    wire n3931 ;
    wire n3932 ;
    wire n3933 ;
    wire n3934 ;
    wire n3935 ;
    wire n3936 ;
    wire n3937 ;
    wire n3938 ;
    wire n3939 ;
    wire n3940 ;
    wire n3941 ;
    wire n3942 ;
    wire n3943 ;
    wire n3944 ;
    wire n3945 ;
    wire n3946 ;
    wire n3947 ;
    wire n3948 ;
    wire n3949 ;
    wire n3950 ;
    wire n3951 ;
    wire n3952 ;
    wire n3953 ;
    wire n3954 ;
    wire n3955 ;
    wire n3956 ;
    wire n3957 ;
    wire n3958 ;
    wire n3959 ;
    wire n3960 ;
    wire n3961 ;
    wire n3962 ;
    wire n3963 ;
    wire n3964 ;
    wire n3965 ;
    wire n3966 ;
    wire n3967 ;
    wire n3968 ;
    wire n3969 ;
    wire n3970 ;
    wire n3971 ;
    wire n3972 ;
    wire n3973 ;
    wire n3974 ;
    wire n3975 ;
    wire n3976 ;
    wire n3977 ;
    wire n3978 ;
    wire n3979 ;
    wire n3980 ;
    wire n3981 ;
    wire n3982 ;
    wire n3983 ;
    wire n3984 ;
    wire n3985 ;
    wire n3986 ;
    wire n3987 ;
    wire n3988 ;
    wire n3989 ;
    wire n3990 ;
    wire n3991 ;
    wire n3992 ;
    wire n3993 ;
    wire n3994 ;
    wire n3995 ;
    wire n3996 ;
    wire n3997 ;
    wire n3998 ;
    wire n3999 ;
    wire n4000 ;
    wire n4001 ;
    wire n4002 ;
    wire n4003 ;
    wire n4004 ;
    wire n4005 ;
    wire n4006 ;
    wire n4007 ;
    wire n4008 ;
    wire n4009 ;
    wire n4010 ;
    wire n4011 ;
    wire n4012 ;
    wire n4013 ;
    wire n4014 ;
    wire n4015 ;
    wire n4016 ;
    wire n4017 ;
    wire n4018 ;
    wire n4019 ;
    wire n4020 ;
    wire n4021 ;
    wire n4022 ;
    wire n4023 ;
    wire n4024 ;
    wire n4025 ;
    wire n4026 ;
    wire n4027 ;
    wire n4028 ;
    wire n4029 ;
    wire n4030 ;
    wire n4031 ;
    wire n4032 ;
    wire n4033 ;
    wire n4034 ;
    wire n4035 ;
    wire n4036 ;
    wire n4037 ;
    wire n4038 ;
    wire n4039 ;
    wire n4040 ;
    wire n4041 ;
    wire n4042 ;
    wire n4043 ;
    wire n4044 ;
    wire n4045 ;
    wire n4046 ;
    wire n4047 ;
    wire n4048 ;
    wire n4049 ;
    wire n4050 ;
    wire n4051 ;
    wire n4052 ;
    wire n4053 ;
    wire n4054 ;
    wire n4055 ;
    wire n4056 ;
    wire n4057 ;
    wire n4058 ;
    wire n4059 ;
    wire n4060 ;
    wire n4061 ;
    wire n4062 ;
    wire n4063 ;
    wire n4064 ;
    wire n4065 ;
    wire n4066 ;
    wire n4067 ;
    wire n4068 ;
    wire n4069 ;
    wire n4070 ;
    wire n4071 ;
    wire n4072 ;
    wire n4073 ;
    wire n4074 ;
    wire n4075 ;
    wire n4076 ;
    wire n4077 ;
    wire n4078 ;
    wire n4079 ;
    wire n4080 ;
    wire n4081 ;
    wire n4082 ;
    wire n4083 ;
    wire n4084 ;
    wire n4085 ;
    wire n4086 ;
    wire n4087 ;
    wire n4088 ;
    wire n4089 ;
    wire n4090 ;
    wire n4091 ;
    wire n4092 ;
    wire n4093 ;
    wire n4094 ;
    wire n4095 ;
    wire n4096 ;
    wire n4097 ;
    wire n4098 ;
    wire n4099 ;
    wire n4100 ;
    wire n4101 ;
    wire n4102 ;
    wire n4103 ;
    wire n4104 ;
    wire n4105 ;
    wire n4106 ;
    wire n4107 ;
    wire n4108 ;
    wire n4109 ;
    wire n4110 ;
    wire n4111 ;
    wire n4112 ;
    wire n4113 ;
    wire n4114 ;
    wire n4115 ;
    wire n4116 ;
    wire n4117 ;
    wire n4118 ;
    wire n4119 ;
    wire n4120 ;
    wire n4121 ;
    wire n4122 ;
    wire n4123 ;
    wire n4124 ;
    wire n4125 ;
    wire n4126 ;
    wire n4127 ;
    wire n4128 ;
    wire n4129 ;
    wire n4130 ;
    wire n4131 ;
    wire n4132 ;
    wire n4133 ;
    wire n4134 ;
    wire n4135 ;
    wire n4136 ;
    wire n4137 ;
    wire n4138 ;
    wire n4139 ;
    wire n4140 ;
    wire n4141 ;
    wire n4142 ;
    wire n4143 ;
    wire n4144 ;
    wire n4145 ;
    wire n4146 ;
    wire n4147 ;
    wire n4148 ;
    wire n4149 ;
    wire n4150 ;
    wire n4151 ;
    wire n4152 ;
    wire n4153 ;
    wire n4154 ;
    wire n4155 ;
    wire n4156 ;
    wire n4157 ;
    wire n4158 ;
    wire n4159 ;
    wire n4160 ;
    wire n4161 ;
    wire n4162 ;
    wire n4163 ;
    wire n4164 ;
    wire n4165 ;
    wire n4166 ;
    wire n4167 ;
    wire n4168 ;
    wire n4169 ;
    wire n4170 ;
    wire n4171 ;
    wire n4172 ;
    wire n4173 ;
    wire n4174 ;
    wire n4175 ;
    wire n4176 ;
    wire n4177 ;
    wire n4178 ;
    wire n4179 ;
    wire n4180 ;
    wire n4181 ;
    wire n4182 ;
    wire n4183 ;
    wire n4184 ;
    wire n4185 ;
    wire n4186 ;
    wire n4187 ;
    wire n4188 ;
    wire n4189 ;
    wire n4190 ;
    wire n4191 ;
    wire n4192 ;
    wire n4193 ;
    wire n4194 ;
    wire n4195 ;
    wire n4196 ;
    wire n4197 ;
    wire n4198 ;
    wire n4199 ;
    wire n4200 ;
    wire n4201 ;
    wire n4202 ;
    wire n4203 ;
    wire n4204 ;
    wire n4205 ;
    wire n4206 ;
    wire n4207 ;
    wire n4208 ;
    wire n4209 ;
    wire n4210 ;
    wire n4211 ;
    wire n4212 ;
    wire n4213 ;
    wire n4214 ;
    wire n4215 ;
    wire n4216 ;
    wire n4217 ;
    wire n4218 ;
    wire n4219 ;
    wire n4220 ;
    wire n4221 ;
    wire n4222 ;
    wire n4223 ;
    wire n4224 ;
    wire n4225 ;
    wire n4226 ;
    wire n4227 ;
    wire n4228 ;
    wire n4229 ;
    wire n4230 ;
    wire n4231 ;
    wire n4232 ;
    wire n4233 ;
    wire n4234 ;
    wire n4235 ;
    wire n4236 ;
    wire n4237 ;
    wire n4238 ;
    wire n4239 ;
    wire n4240 ;
    wire n4241 ;
    wire n4242 ;
    wire n4243 ;
    wire n4244 ;
    wire n4245 ;
    wire n4246 ;
    wire n4247 ;
    wire n4248 ;
    wire n4249 ;
    wire n4250 ;
    wire n4251 ;
    wire n4252 ;
    wire n4253 ;
    wire n4254 ;
    wire n4255 ;
    wire n4256 ;
    wire n4257 ;
    wire n4258 ;
    wire n4259 ;
    wire n4260 ;
    wire n4261 ;
    wire n4262 ;
    wire n4263 ;
    wire n4264 ;
    wire n4265 ;
    wire n4266 ;
    wire n4267 ;
    wire n4268 ;
    wire n4269 ;
    wire n4270 ;
    wire n4271 ;
    wire n4272 ;
    wire SboxInst_n384 ;
    wire SboxInst_n383 ;
    wire SboxInst_n382 ;
    wire SboxInst_n381 ;
    wire SboxInst_n380 ;
    wire SboxInst_n379 ;
    wire SboxInst_n378 ;
    wire SboxInst_n377 ;
    wire SboxInst_n376 ;
    wire SboxInst_n375 ;
    wire SboxInst_n374 ;
    wire SboxInst_n373 ;
    wire SboxInst_n372 ;
    wire SboxInst_n371 ;
    wire SboxInst_n370 ;
    wire SboxInst_n369 ;
    wire SboxInst_n368 ;
    wire SboxInst_n367 ;
    wire SboxInst_n366 ;
    wire SboxInst_n365 ;
    wire SboxInst_n364 ;
    wire SboxInst_n363 ;
    wire SboxInst_n362 ;
    wire SboxInst_n361 ;
    wire SboxInst_n360 ;
    wire SboxInst_n359 ;
    wire SboxInst_n358 ;
    wire SboxInst_n357 ;
    wire SboxInst_n356 ;
    wire SboxInst_n355 ;
    wire SboxInst_n354 ;
    wire SboxInst_n353 ;
    wire SboxInst_n352 ;
    wire SboxInst_n351 ;
    wire SboxInst_n350 ;
    wire SboxInst_n349 ;
    wire SboxInst_n348 ;
    wire SboxInst_n347 ;
    wire SboxInst_n346 ;
    wire SboxInst_n345 ;
    wire SboxInst_n344 ;
    wire SboxInst_n343 ;
    wire SboxInst_n342 ;
    wire SboxInst_n341 ;
    wire SboxInst_n340 ;
    wire SboxInst_n339 ;
    wire SboxInst_n338 ;
    wire SboxInst_n337 ;
    wire SboxInst_n336 ;
    wire SboxInst_n335 ;
    wire SboxInst_n334 ;
    wire SboxInst_n333 ;
    wire SboxInst_n332 ;
    wire SboxInst_n331 ;
    wire SboxInst_n330 ;
    wire SboxInst_n329 ;
    wire SboxInst_n328 ;
    wire SboxInst_n327 ;
    wire SboxInst_n326 ;
    wire SboxInst_n325 ;
    wire SboxInst_n324 ;
    wire SboxInst_n323 ;
    wire SboxInst_n322 ;
    wire SboxInst_n321 ;
    wire SboxInst_n320 ;
    wire SboxInst_n319 ;
    wire SboxInst_n318 ;
    wire SboxInst_n317 ;
    wire SboxInst_n316 ;
    wire SboxInst_n315 ;
    wire SboxInst_n314 ;
    wire SboxInst_n313 ;
    wire SboxInst_n312 ;
    wire SboxInst_n311 ;
    wire SboxInst_n310 ;
    wire SboxInst_n309 ;
    wire SboxInst_n308 ;
    wire SboxInst_n307 ;
    wire SboxInst_n306 ;
    wire SboxInst_n305 ;
    wire SboxInst_n304 ;
    wire SboxInst_n303 ;
    wire SboxInst_n302 ;
    wire SboxInst_n301 ;
    wire SboxInst_n300 ;
    wire SboxInst_n299 ;
    wire SboxInst_n298 ;
    wire SboxInst_n297 ;
    wire SboxInst_n296 ;
    wire SboxInst_n295 ;
    wire SboxInst_n294 ;
    wire SboxInst_n293 ;
    wire SboxInst_n292 ;
    wire SboxInst_n291 ;
    wire SboxInst_n290 ;
    wire SboxInst_n289 ;
    wire SboxInst_n288 ;
    wire SboxInst_n287 ;
    wire SboxInst_n286 ;
    wire SboxInst_n285 ;
    wire SboxInst_n284 ;
    wire SboxInst_n283 ;
    wire SboxInst_n282 ;
    wire SboxInst_n281 ;
    wire SboxInst_n280 ;
    wire SboxInst_n279 ;
    wire SboxInst_n278 ;
    wire SboxInst_n277 ;
    wire SboxInst_n276 ;
    wire SboxInst_n275 ;
    wire SboxInst_n274 ;
    wire SboxInst_n273 ;
    wire SboxInst_n272 ;
    wire SboxInst_n271 ;
    wire SboxInst_n270 ;
    wire SboxInst_n269 ;
    wire SboxInst_n268 ;
    wire SboxInst_n267 ;
    wire SboxInst_n266 ;
    wire SboxInst_n265 ;
    wire SboxInst_n264 ;
    wire SboxInst_n263 ;
    wire SboxInst_n262 ;
    wire SboxInst_n261 ;
    wire SboxInst_n260 ;
    wire SboxInst_n259 ;
    wire SboxInst_n258 ;
    wire SboxInst_n257 ;
    wire SboxInst_n256 ;
    wire SboxInst_n255 ;
    wire SboxInst_n254 ;
    wire SboxInst_n253 ;
    wire SboxInst_n252 ;
    wire SboxInst_n251 ;
    wire SboxInst_n250 ;
    wire SboxInst_n249 ;
    wire SboxInst_n248 ;
    wire SboxInst_n247 ;
    wire SboxInst_n246 ;
    wire SboxInst_n245 ;
    wire SboxInst_n244 ;
    wire SboxInst_n243 ;
    wire SboxInst_n242 ;
    wire SboxInst_n241 ;
    wire SboxInst_n240 ;
    wire SboxInst_n239 ;
    wire SboxInst_n238 ;
    wire SboxInst_n237 ;
    wire SboxInst_n236 ;
    wire SboxInst_n235 ;
    wire SboxInst_n234 ;
    wire SboxInst_n233 ;
    wire SboxInst_n232 ;
    wire SboxInst_n231 ;
    wire SboxInst_n230 ;
    wire SboxInst_n229 ;
    wire SboxInst_n228 ;
    wire SboxInst_n227 ;
    wire SboxInst_n226 ;
    wire SboxInst_n225 ;
    wire SboxInst_n224 ;
    wire SboxInst_n223 ;
    wire SboxInst_n222 ;
    wire SboxInst_n221 ;
    wire SboxInst_n220 ;
    wire SboxInst_n219 ;
    wire SboxInst_n218 ;
    wire SboxInst_n217 ;
    wire SboxInst_n216 ;
    wire SboxInst_n215 ;
    wire SboxInst_n214 ;
    wire SboxInst_n213 ;
    wire SboxInst_n212 ;
    wire SboxInst_n211 ;
    wire SboxInst_n210 ;
    wire SboxInst_n209 ;
    wire SboxInst_n208 ;
    wire SboxInst_n207 ;
    wire SboxInst_n206 ;
    wire SboxInst_n205 ;
    wire SboxInst_n204 ;
    wire SboxInst_n203 ;
    wire SboxInst_n202 ;
    wire SboxInst_n201 ;
    wire SboxInst_n200 ;
    wire SboxInst_n199 ;
    wire SboxInst_n198 ;
    wire SboxInst_n197 ;
    wire SboxInst_n196 ;
    wire SboxInst_n195 ;
    wire SboxInst_n194 ;
    wire SboxInst_n193 ;
    wire [63:0] y0 ;
    wire [1:0] y2 ;
    wire [63:0] y4 ;
    wire [63:0] z0 ;
    wire [63:0] z1 ;
    wire [63:0] z2 ;
    wire [63:0] z3 ;
    wire [63:0] z4 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4651 ;
    wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 U3097 ( .a ({state_in_s1[241], state_in_s0[241]}), .b ({state_in_s1[305], state_in_s0[305]}), .c ({new_AGEMA_signal_2338, y4[9]}) ) ;
    xor_HPC2 U3098 ( .a ({state_in_s1[304], state_in_s0[304]}), .b ({state_in_s1[240], state_in_s0[240]}), .c ({new_AGEMA_signal_2341, y4[8]}) ) ;
    xor_HPC2 U3099 ( .a ({state_in_s1[255], state_in_s0[255]}), .b ({state_in_s1[319], state_in_s0[319]}), .c ({new_AGEMA_signal_2344, y4[7]}) ) ;
    xor_HPC2 U3100 ( .a ({state_in_s1[254], state_in_s0[254]}), .b ({state_in_s1[318], state_in_s0[318]}), .c ({new_AGEMA_signal_2347, y4[6]}) ) ;
    xor_HPC2 U3101 ( .a ({state_in_s1[199], state_in_s0[199]}), .b ({state_in_s1[263], state_in_s0[263]}), .c ({new_AGEMA_signal_2350, y4[63]}) ) ;
    xor_HPC2 U3102 ( .a ({state_in_s1[262], state_in_s0[262]}), .b ({state_in_s1[198], state_in_s0[198]}), .c ({new_AGEMA_signal_2353, y4[62]}) ) ;
    xor_HPC2 U3103 ( .a ({state_in_s1[197], state_in_s0[197]}), .b ({state_in_s1[261], state_in_s0[261]}), .c ({new_AGEMA_signal_2356, y4[61]}) ) ;
    xor_HPC2 U3104 ( .a ({state_in_s1[196], state_in_s0[196]}), .b ({state_in_s1[260], state_in_s0[260]}), .c ({new_AGEMA_signal_2359, y4[60]}) ) ;
    xor_HPC2 U3105 ( .a ({state_in_s1[317], state_in_s0[317]}), .b ({state_in_s1[253], state_in_s0[253]}), .c ({new_AGEMA_signal_2362, y4[5]}) ) ;
    xor_HPC2 U3106 ( .a ({state_in_s1[195], state_in_s0[195]}), .b ({state_in_s1[259], state_in_s0[259]}), .c ({new_AGEMA_signal_2365, y4[59]}) ) ;
    xor_HPC2 U3107 ( .a ({state_in_s1[258], state_in_s0[258]}), .b ({state_in_s1[194], state_in_s0[194]}), .c ({new_AGEMA_signal_2368, y4[58]}) ) ;
    xor_HPC2 U3108 ( .a ({state_in_s1[193], state_in_s0[193]}), .b ({state_in_s1[257], state_in_s0[257]}), .c ({new_AGEMA_signal_2371, y4[57]}) ) ;
    xor_HPC2 U3109 ( .a ({state_in_s1[192], state_in_s0[192]}), .b ({state_in_s1[256], state_in_s0[256]}), .c ({new_AGEMA_signal_2374, y4[56]}) ) ;
    xor_HPC2 U3110 ( .a ({state_in_s1[271], state_in_s0[271]}), .b ({state_in_s1[207], state_in_s0[207]}), .c ({new_AGEMA_signal_2377, y4[55]}) ) ;
    xor_HPC2 U3111 ( .a ({state_in_s1[206], state_in_s0[206]}), .b ({state_in_s1[270], state_in_s0[270]}), .c ({new_AGEMA_signal_2380, y4[54]}) ) ;
    xor_HPC2 U3112 ( .a ({state_in_s1[205], state_in_s0[205]}), .b ({state_in_s1[269], state_in_s0[269]}), .c ({new_AGEMA_signal_2383, y4[53]}) ) ;
    xor_HPC2 U3113 ( .a ({state_in_s1[268], state_in_s0[268]}), .b ({state_in_s1[204], state_in_s0[204]}), .c ({new_AGEMA_signal_2386, y4[52]}) ) ;
    xor_HPC2 U3114 ( .a ({state_in_s1[267], state_in_s0[267]}), .b ({state_in_s1[203], state_in_s0[203]}), .c ({new_AGEMA_signal_2389, y4[51]}) ) ;
    xor_HPC2 U3115 ( .a ({state_in_s1[202], state_in_s0[202]}), .b ({state_in_s1[266], state_in_s0[266]}), .c ({new_AGEMA_signal_2392, y4[50]}) ) ;
    xor_HPC2 U3116 ( .a ({state_in_s1[316], state_in_s0[316]}), .b ({state_in_s1[252], state_in_s0[252]}), .c ({new_AGEMA_signal_2395, y4[4]}) ) ;
    xor_HPC2 U3117 ( .a ({state_in_s1[201], state_in_s0[201]}), .b ({state_in_s1[265], state_in_s0[265]}), .c ({new_AGEMA_signal_2398, y4[49]}) ) ;
    xor_HPC2 U3118 ( .a ({state_in_s1[264], state_in_s0[264]}), .b ({state_in_s1[200], state_in_s0[200]}), .c ({new_AGEMA_signal_2401, y4[48]}) ) ;
    xor_HPC2 U3119 ( .a ({state_in_s1[279], state_in_s0[279]}), .b ({state_in_s1[215], state_in_s0[215]}), .c ({new_AGEMA_signal_2404, y4[47]}) ) ;
    xor_HPC2 U3120 ( .a ({state_in_s1[278], state_in_s0[278]}), .b ({state_in_s1[214], state_in_s0[214]}), .c ({new_AGEMA_signal_2407, y4[46]}) ) ;
    xor_HPC2 U3121 ( .a ({state_in_s1[277], state_in_s0[277]}), .b ({state_in_s1[213], state_in_s0[213]}), .c ({new_AGEMA_signal_2410, y4[45]}) ) ;
    xor_HPC2 U3122 ( .a ({state_in_s1[276], state_in_s0[276]}), .b ({state_in_s1[212], state_in_s0[212]}), .c ({new_AGEMA_signal_2413, y4[44]}) ) ;
    xor_HPC2 U3123 ( .a ({state_in_s1[275], state_in_s0[275]}), .b ({state_in_s1[211], state_in_s0[211]}), .c ({new_AGEMA_signal_2416, y4[43]}) ) ;
    xor_HPC2 U3124 ( .a ({state_in_s1[274], state_in_s0[274]}), .b ({state_in_s1[210], state_in_s0[210]}), .c ({new_AGEMA_signal_2419, y4[42]}) ) ;
    xor_HPC2 U3125 ( .a ({state_in_s1[273], state_in_s0[273]}), .b ({state_in_s1[209], state_in_s0[209]}), .c ({new_AGEMA_signal_2422, y4[41]}) ) ;
    xor_HPC2 U3126 ( .a ({state_in_s1[272], state_in_s0[272]}), .b ({state_in_s1[208], state_in_s0[208]}), .c ({new_AGEMA_signal_2425, y4[40]}) ) ;
    xor_HPC2 U3127 ( .a ({state_in_s1[251], state_in_s0[251]}), .b ({state_in_s1[315], state_in_s0[315]}), .c ({new_AGEMA_signal_2428, y4[3]}) ) ;
    xor_HPC2 U3128 ( .a ({state_in_s1[287], state_in_s0[287]}), .b ({state_in_s1[223], state_in_s0[223]}), .c ({new_AGEMA_signal_2431, y4[39]}) ) ;
    xor_HPC2 U3129 ( .a ({state_in_s1[286], state_in_s0[286]}), .b ({state_in_s1[222], state_in_s0[222]}), .c ({new_AGEMA_signal_2434, y4[38]}) ) ;
    xor_HPC2 U3130 ( .a ({state_in_s1[285], state_in_s0[285]}), .b ({state_in_s1[221], state_in_s0[221]}), .c ({new_AGEMA_signal_2437, y4[37]}) ) ;
    xor_HPC2 U3131 ( .a ({state_in_s1[284], state_in_s0[284]}), .b ({state_in_s1[220], state_in_s0[220]}), .c ({new_AGEMA_signal_2440, y4[36]}) ) ;
    xor_HPC2 U3132 ( .a ({state_in_s1[283], state_in_s0[283]}), .b ({state_in_s1[219], state_in_s0[219]}), .c ({new_AGEMA_signal_2443, y4[35]}) ) ;
    xor_HPC2 U3133 ( .a ({state_in_s1[282], state_in_s0[282]}), .b ({state_in_s1[218], state_in_s0[218]}), .c ({new_AGEMA_signal_2446, y4[34]}) ) ;
    xor_HPC2 U3134 ( .a ({state_in_s1[281], state_in_s0[281]}), .b ({state_in_s1[217], state_in_s0[217]}), .c ({new_AGEMA_signal_2449, y4[33]}) ) ;
    xor_HPC2 U3135 ( .a ({state_in_s1[280], state_in_s0[280]}), .b ({state_in_s1[216], state_in_s0[216]}), .c ({new_AGEMA_signal_2452, y4[32]}) ) ;
    xor_HPC2 U3136 ( .a ({state_in_s1[295], state_in_s0[295]}), .b ({state_in_s1[231], state_in_s0[231]}), .c ({new_AGEMA_signal_2455, y4[31]}) ) ;
    xor_HPC2 U3137 ( .a ({state_in_s1[294], state_in_s0[294]}), .b ({state_in_s1[230], state_in_s0[230]}), .c ({new_AGEMA_signal_2458, y4[30]}) ) ;
    xor_HPC2 U3138 ( .a ({state_in_s1[250], state_in_s0[250]}), .b ({state_in_s1[314], state_in_s0[314]}), .c ({new_AGEMA_signal_2461, y4[2]}) ) ;
    xor_HPC2 U3139 ( .a ({state_in_s1[293], state_in_s0[293]}), .b ({state_in_s1[229], state_in_s0[229]}), .c ({new_AGEMA_signal_2464, y4[29]}) ) ;
    xor_HPC2 U3140 ( .a ({state_in_s1[292], state_in_s0[292]}), .b ({state_in_s1[228], state_in_s0[228]}), .c ({new_AGEMA_signal_2467, y4[28]}) ) ;
    xor_HPC2 U3141 ( .a ({state_in_s1[291], state_in_s0[291]}), .b ({state_in_s1[227], state_in_s0[227]}), .c ({new_AGEMA_signal_2470, y4[27]}) ) ;
    xor_HPC2 U3142 ( .a ({state_in_s1[290], state_in_s0[290]}), .b ({state_in_s1[226], state_in_s0[226]}), .c ({new_AGEMA_signal_2473, y4[26]}) ) ;
    xor_HPC2 U3143 ( .a ({state_in_s1[289], state_in_s0[289]}), .b ({state_in_s1[225], state_in_s0[225]}), .c ({new_AGEMA_signal_2476, y4[25]}) ) ;
    xor_HPC2 U3144 ( .a ({state_in_s1[224], state_in_s0[224]}), .b ({state_in_s1[288], state_in_s0[288]}), .c ({new_AGEMA_signal_2479, y4[24]}) ) ;
    xor_HPC2 U3145 ( .a ({state_in_s1[239], state_in_s0[239]}), .b ({state_in_s1[303], state_in_s0[303]}), .c ({new_AGEMA_signal_2482, y4[23]}) ) ;
    xor_HPC2 U3146 ( .a ({state_in_s1[302], state_in_s0[302]}), .b ({state_in_s1[238], state_in_s0[238]}), .c ({new_AGEMA_signal_2485, y4[22]}) ) ;
    xor_HPC2 U3147 ( .a ({state_in_s1[301], state_in_s0[301]}), .b ({state_in_s1[237], state_in_s0[237]}), .c ({new_AGEMA_signal_2488, y4[21]}) ) ;
    xor_HPC2 U3148 ( .a ({state_in_s1[236], state_in_s0[236]}), .b ({state_in_s1[300], state_in_s0[300]}), .c ({new_AGEMA_signal_2491, y4[20]}) ) ;
    xor_HPC2 U3149 ( .a ({state_in_s1[313], state_in_s0[313]}), .b ({state_in_s1[249], state_in_s0[249]}), .c ({new_AGEMA_signal_2494, y4[1]}) ) ;
    xor_HPC2 U3150 ( .a ({state_in_s1[235], state_in_s0[235]}), .b ({state_in_s1[299], state_in_s0[299]}), .c ({new_AGEMA_signal_2497, y4[19]}) ) ;
    xor_HPC2 U3151 ( .a ({state_in_s1[298], state_in_s0[298]}), .b ({state_in_s1[234], state_in_s0[234]}), .c ({new_AGEMA_signal_2500, y4[18]}) ) ;
    xor_HPC2 U3152 ( .a ({state_in_s1[233], state_in_s0[233]}), .b ({state_in_s1[297], state_in_s0[297]}), .c ({new_AGEMA_signal_2503, y4[17]}) ) ;
    xor_HPC2 U3153 ( .a ({state_in_s1[232], state_in_s0[232]}), .b ({state_in_s1[296], state_in_s0[296]}), .c ({new_AGEMA_signal_2506, y4[16]}) ) ;
    xor_HPC2 U3154 ( .a ({state_in_s1[311], state_in_s0[311]}), .b ({state_in_s1[247], state_in_s0[247]}), .c ({new_AGEMA_signal_2509, y4[15]}) ) ;
    xor_HPC2 U3155 ( .a ({state_in_s1[246], state_in_s0[246]}), .b ({state_in_s1[310], state_in_s0[310]}), .c ({new_AGEMA_signal_2512, y4[14]}) ) ;
    xor_HPC2 U3156 ( .a ({state_in_s1[245], state_in_s0[245]}), .b ({state_in_s1[309], state_in_s0[309]}), .c ({new_AGEMA_signal_2515, y4[13]}) ) ;
    xor_HPC2 U3157 ( .a ({state_in_s1[244], state_in_s0[244]}), .b ({state_in_s1[308], state_in_s0[308]}), .c ({new_AGEMA_signal_2518, y4[12]}) ) ;
    xor_HPC2 U3158 ( .a ({state_in_s1[307], state_in_s0[307]}), .b ({state_in_s1[243], state_in_s0[243]}), .c ({new_AGEMA_signal_2521, y4[11]}) ) ;
    xor_HPC2 U3159 ( .a ({state_in_s1[242], state_in_s0[242]}), .b ({state_in_s1[306], state_in_s0[306]}), .c ({new_AGEMA_signal_2524, y4[10]}) ) ;
    xor_HPC2 U3160 ( .a ({state_in_s1[248], state_in_s0[248]}), .b ({state_in_s1[312], state_in_s0[312]}), .c ({new_AGEMA_signal_2527, y4[0]}) ) ;
    xor_HPC2 U3161 ( .a ({state_in_s1[49], state_in_s0[49]}), .b ({state_in_s1[305], state_in_s0[305]}), .c ({new_AGEMA_signal_2529, y0[9]}) ) ;
    xor_HPC2 U3162 ( .a ({state_in_s1[48], state_in_s0[48]}), .b ({state_in_s1[304], state_in_s0[304]}), .c ({new_AGEMA_signal_2531, y0[8]}) ) ;
    xor_HPC2 U3163 ( .a ({state_in_s1[63], state_in_s0[63]}), .b ({state_in_s1[319], state_in_s0[319]}), .c ({new_AGEMA_signal_2533, y0[7]}) ) ;
    xor_HPC2 U3164 ( .a ({state_in_s1[62], state_in_s0[62]}), .b ({state_in_s1[318], state_in_s0[318]}), .c ({new_AGEMA_signal_2535, y0[6]}) ) ;
    xor_HPC2 U3165 ( .a ({state_in_s1[7], state_in_s0[7]}), .b ({state_in_s1[263], state_in_s0[263]}), .c ({new_AGEMA_signal_2537, y0[63]}) ) ;
    xor_HPC2 U3166 ( .a ({state_in_s1[6], state_in_s0[6]}), .b ({state_in_s1[262], state_in_s0[262]}), .c ({new_AGEMA_signal_2539, y0[62]}) ) ;
    xor_HPC2 U3167 ( .a ({state_in_s1[5], state_in_s0[5]}), .b ({state_in_s1[261], state_in_s0[261]}), .c ({new_AGEMA_signal_2541, y0[61]}) ) ;
    xor_HPC2 U3168 ( .a ({state_in_s1[4], state_in_s0[4]}), .b ({state_in_s1[260], state_in_s0[260]}), .c ({new_AGEMA_signal_2543, y0[60]}) ) ;
    xor_HPC2 U3169 ( .a ({state_in_s1[61], state_in_s0[61]}), .b ({state_in_s1[317], state_in_s0[317]}), .c ({new_AGEMA_signal_2545, y0[5]}) ) ;
    xor_HPC2 U3170 ( .a ({state_in_s1[259], state_in_s0[259]}), .b ({state_in_s1[3], state_in_s0[3]}), .c ({new_AGEMA_signal_2547, y0[59]}) ) ;
    xor_HPC2 U3171 ( .a ({state_in_s1[258], state_in_s0[258]}), .b ({state_in_s1[2], state_in_s0[2]}), .c ({new_AGEMA_signal_2549, y0[58]}) ) ;
    xor_HPC2 U3172 ( .a ({state_in_s1[257], state_in_s0[257]}), .b ({state_in_s1[1], state_in_s0[1]}), .c ({new_AGEMA_signal_2551, y0[57]}) ) ;
    xor_HPC2 U3173 ( .a ({state_in_s1[0], state_in_s0[0]}), .b ({state_in_s1[256], state_in_s0[256]}), .c ({new_AGEMA_signal_2553, y0[56]}) ) ;
    xor_HPC2 U3174 ( .a ({state_in_s1[15], state_in_s0[15]}), .b ({state_in_s1[271], state_in_s0[271]}), .c ({new_AGEMA_signal_2555, y0[55]}) ) ;
    xor_HPC2 U3175 ( .a ({state_in_s1[14], state_in_s0[14]}), .b ({state_in_s1[270], state_in_s0[270]}), .c ({new_AGEMA_signal_2557, y0[54]}) ) ;
    xor_HPC2 U3176 ( .a ({state_in_s1[13], state_in_s0[13]}), .b ({state_in_s1[269], state_in_s0[269]}), .c ({new_AGEMA_signal_2559, y0[53]}) ) ;
    xor_HPC2 U3177 ( .a ({state_in_s1[268], state_in_s0[268]}), .b ({state_in_s1[12], state_in_s0[12]}), .c ({new_AGEMA_signal_2561, y0[52]}) ) ;
    xor_HPC2 U3178 ( .a ({state_in_s1[267], state_in_s0[267]}), .b ({state_in_s1[11], state_in_s0[11]}), .c ({new_AGEMA_signal_2563, y0[51]}) ) ;
    xor_HPC2 U3179 ( .a ({state_in_s1[10], state_in_s0[10]}), .b ({state_in_s1[266], state_in_s0[266]}), .c ({new_AGEMA_signal_2565, y0[50]}) ) ;
    xor_HPC2 U3180 ( .a ({state_in_s1[60], state_in_s0[60]}), .b ({state_in_s1[316], state_in_s0[316]}), .c ({new_AGEMA_signal_2567, y0[4]}) ) ;
    xor_HPC2 U3181 ( .a ({state_in_s1[9], state_in_s0[9]}), .b ({state_in_s1[265], state_in_s0[265]}), .c ({new_AGEMA_signal_2569, y0[49]}) ) ;
    xor_HPC2 U3182 ( .a ({state_in_s1[264], state_in_s0[264]}), .b ({state_in_s1[8], state_in_s0[8]}), .c ({new_AGEMA_signal_2571, y0[48]}) ) ;
    xor_HPC2 U3183 ( .a ({state_in_s1[279], state_in_s0[279]}), .b ({state_in_s1[23], state_in_s0[23]}), .c ({new_AGEMA_signal_2573, y0[47]}) ) ;
    xor_HPC2 U3184 ( .a ({state_in_s1[22], state_in_s0[22]}), .b ({state_in_s1[278], state_in_s0[278]}), .c ({new_AGEMA_signal_2575, y0[46]}) ) ;
    xor_HPC2 U3185 ( .a ({state_in_s1[277], state_in_s0[277]}), .b ({state_in_s1[21], state_in_s0[21]}), .c ({new_AGEMA_signal_2577, y0[45]}) ) ;
    xor_HPC2 U3186 ( .a ({state_in_s1[276], state_in_s0[276]}), .b ({state_in_s1[20], state_in_s0[20]}), .c ({new_AGEMA_signal_2579, y0[44]}) ) ;
    xor_HPC2 U3187 ( .a ({state_in_s1[19], state_in_s0[19]}), .b ({state_in_s1[275], state_in_s0[275]}), .c ({new_AGEMA_signal_2581, y0[43]}) ) ;
    xor_HPC2 U3188 ( .a ({state_in_s1[18], state_in_s0[18]}), .b ({state_in_s1[274], state_in_s0[274]}), .c ({new_AGEMA_signal_2583, y0[42]}) ) ;
    xor_HPC2 U3189 ( .a ({state_in_s1[273], state_in_s0[273]}), .b ({state_in_s1[17], state_in_s0[17]}), .c ({new_AGEMA_signal_2585, y0[41]}) ) ;
    xor_HPC2 U3190 ( .a ({state_in_s1[16], state_in_s0[16]}), .b ({state_in_s1[272], state_in_s0[272]}), .c ({new_AGEMA_signal_2587, y0[40]}) ) ;
    xor_HPC2 U3191 ( .a ({state_in_s1[59], state_in_s0[59]}), .b ({state_in_s1[315], state_in_s0[315]}), .c ({new_AGEMA_signal_2589, y0[3]}) ) ;
    xor_HPC2 U3192 ( .a ({state_in_s1[31], state_in_s0[31]}), .b ({state_in_s1[287], state_in_s0[287]}), .c ({new_AGEMA_signal_2591, y0[39]}) ) ;
    xor_HPC2 U3193 ( .a ({state_in_s1[30], state_in_s0[30]}), .b ({state_in_s1[286], state_in_s0[286]}), .c ({new_AGEMA_signal_2593, y0[38]}) ) ;
    xor_HPC2 U3194 ( .a ({state_in_s1[29], state_in_s0[29]}), .b ({state_in_s1[285], state_in_s0[285]}), .c ({new_AGEMA_signal_2595, y0[37]}) ) ;
    xor_HPC2 U3195 ( .a ({state_in_s1[28], state_in_s0[28]}), .b ({state_in_s1[284], state_in_s0[284]}), .c ({new_AGEMA_signal_2597, y0[36]}) ) ;
    xor_HPC2 U3196 ( .a ({state_in_s1[27], state_in_s0[27]}), .b ({state_in_s1[283], state_in_s0[283]}), .c ({new_AGEMA_signal_2599, y0[35]}) ) ;
    xor_HPC2 U3197 ( .a ({state_in_s1[26], state_in_s0[26]}), .b ({state_in_s1[282], state_in_s0[282]}), .c ({new_AGEMA_signal_2601, y0[34]}) ) ;
    xor_HPC2 U3198 ( .a ({state_in_s1[25], state_in_s0[25]}), .b ({state_in_s1[281], state_in_s0[281]}), .c ({new_AGEMA_signal_2603, y0[33]}) ) ;
    xor_HPC2 U3199 ( .a ({state_in_s1[24], state_in_s0[24]}), .b ({state_in_s1[280], state_in_s0[280]}), .c ({new_AGEMA_signal_2605, y0[32]}) ) ;
    xor_HPC2 U3200 ( .a ({state_in_s1[39], state_in_s0[39]}), .b ({state_in_s1[295], state_in_s0[295]}), .c ({new_AGEMA_signal_2607, y0[31]}) ) ;
    xor_HPC2 U3201 ( .a ({state_in_s1[38], state_in_s0[38]}), .b ({state_in_s1[294], state_in_s0[294]}), .c ({new_AGEMA_signal_2609, y0[30]}) ) ;
    xor_HPC2 U3202 ( .a ({state_in_s1[58], state_in_s0[58]}), .b ({state_in_s1[314], state_in_s0[314]}), .c ({new_AGEMA_signal_2611, y0[2]}) ) ;
    xor_HPC2 U3203 ( .a ({state_in_s1[293], state_in_s0[293]}), .b ({state_in_s1[37], state_in_s0[37]}), .c ({new_AGEMA_signal_2613, y0[29]}) ) ;
    xor_HPC2 U3204 ( .a ({state_in_s1[292], state_in_s0[292]}), .b ({state_in_s1[36], state_in_s0[36]}), .c ({new_AGEMA_signal_2615, y0[28]}) ) ;
    xor_HPC2 U3205 ( .a ({state_in_s1[35], state_in_s0[35]}), .b ({state_in_s1[291], state_in_s0[291]}), .c ({new_AGEMA_signal_2617, y0[27]}) ) ;
    xor_HPC2 U3206 ( .a ({state_in_s1[34], state_in_s0[34]}), .b ({state_in_s1[290], state_in_s0[290]}), .c ({new_AGEMA_signal_2619, y0[26]}) ) ;
    xor_HPC2 U3207 ( .a ({state_in_s1[289], state_in_s0[289]}), .b ({state_in_s1[33], state_in_s0[33]}), .c ({new_AGEMA_signal_2621, y0[25]}) ) ;
    xor_HPC2 U3208 ( .a ({state_in_s1[32], state_in_s0[32]}), .b ({state_in_s1[288], state_in_s0[288]}), .c ({new_AGEMA_signal_2623, y0[24]}) ) ;
    xor_HPC2 U3209 ( .a ({state_in_s1[47], state_in_s0[47]}), .b ({state_in_s1[303], state_in_s0[303]}), .c ({new_AGEMA_signal_2625, y0[23]}) ) ;
    xor_HPC2 U3210 ( .a ({state_in_s1[302], state_in_s0[302]}), .b ({state_in_s1[46], state_in_s0[46]}), .c ({new_AGEMA_signal_2627, y0[22]}) ) ;
    xor_HPC2 U3211 ( .a ({state_in_s1[45], state_in_s0[45]}), .b ({state_in_s1[301], state_in_s0[301]}), .c ({new_AGEMA_signal_2629, y0[21]}) ) ;
    xor_HPC2 U3212 ( .a ({state_in_s1[44], state_in_s0[44]}), .b ({state_in_s1[300], state_in_s0[300]}), .c ({new_AGEMA_signal_2631, y0[20]}) ) ;
    xor_HPC2 U3213 ( .a ({state_in_s1[57], state_in_s0[57]}), .b ({state_in_s1[313], state_in_s0[313]}), .c ({new_AGEMA_signal_2633, y0[1]}) ) ;
    xor_HPC2 U3214 ( .a ({state_in_s1[43], state_in_s0[43]}), .b ({state_in_s1[299], state_in_s0[299]}), .c ({new_AGEMA_signal_2635, y0[19]}) ) ;
    xor_HPC2 U3215 ( .a ({state_in_s1[298], state_in_s0[298]}), .b ({state_in_s1[42], state_in_s0[42]}), .c ({new_AGEMA_signal_2637, y0[18]}) ) ;
    xor_HPC2 U3216 ( .a ({state_in_s1[297], state_in_s0[297]}), .b ({state_in_s1[41], state_in_s0[41]}), .c ({new_AGEMA_signal_2639, y0[17]}) ) ;
    xor_HPC2 U3217 ( .a ({state_in_s1[40], state_in_s0[40]}), .b ({state_in_s1[296], state_in_s0[296]}), .c ({new_AGEMA_signal_2641, y0[16]}) ) ;
    xor_HPC2 U3218 ( .a ({state_in_s1[55], state_in_s0[55]}), .b ({state_in_s1[311], state_in_s0[311]}), .c ({new_AGEMA_signal_2643, y0[15]}) ) ;
    xor_HPC2 U3219 ( .a ({state_in_s1[54], state_in_s0[54]}), .b ({state_in_s1[310], state_in_s0[310]}), .c ({new_AGEMA_signal_2645, y0[14]}) ) ;
    xor_HPC2 U3220 ( .a ({state_in_s1[53], state_in_s0[53]}), .b ({state_in_s1[309], state_in_s0[309]}), .c ({new_AGEMA_signal_2647, y0[13]}) ) ;
    xor_HPC2 U3221 ( .a ({state_in_s1[52], state_in_s0[52]}), .b ({state_in_s1[308], state_in_s0[308]}), .c ({new_AGEMA_signal_2649, y0[12]}) ) ;
    xor_HPC2 U3222 ( .a ({state_in_s1[307], state_in_s0[307]}), .b ({state_in_s1[51], state_in_s0[51]}), .c ({new_AGEMA_signal_2651, y0[11]}) ) ;
    xor_HPC2 U3223 ( .a ({state_in_s1[50], state_in_s0[50]}), .b ({state_in_s1[306], state_in_s0[306]}), .c ({new_AGEMA_signal_2653, y0[10]}) ) ;
    xor_HPC2 U3224 ( .a ({state_in_s1[56], state_in_s0[56]}), .b ({state_in_s1[312], state_in_s0[312]}), .c ({new_AGEMA_signal_2655, y0[0]}) ) ;
    xnor_HPC2 U3333 ( .a ({state_in_s1[66], state_in_s0[66]}), .b ({state_in_s1[258], state_in_s0[258]}), .c ({new_AGEMA_signal_2657, n3310}) ) ;
    xnor_HPC2 U3347 ( .a ({state_in_s1[67], state_in_s0[67]}), .b ({state_in_s1[259], state_in_s0[259]}), .c ({new_AGEMA_signal_2659, n3317}) ) ;
    xnor_HPC2 U3379 ( .a ({state_in_s1[65], state_in_s0[65]}), .b ({state_in_s1[257], state_in_s0[257]}), .c ({new_AGEMA_signal_2661, n3329}) ) ;
    xnor_HPC2 U3394 ( .a ({state_in_s1[106], state_in_s0[106]}), .b ({state_in_s1[298], state_in_s0[298]}), .c ({new_AGEMA_signal_2663, n3336}) ) ;
    xnor_HPC2 U3420 ( .a ({state_in_s1[105], state_in_s0[105]}), .b ({state_in_s1[297], state_in_s0[297]}), .c ({new_AGEMA_signal_2665, n3348}) ) ;
    xnor_HPC2 U3458 ( .a ({state_in_s1[97], state_in_s0[97]}), .b ({state_in_s1[289], state_in_s0[289]}), .c ({new_AGEMA_signal_2667, n3367}) ) ;
    xnor_HPC2 U3461 ( .a ({state_in_s1[87], state_in_s0[87]}), .b ({state_in_s1[279], state_in_s0[279]}), .c ({new_AGEMA_signal_2669, n3370}) ) ;
    xnor_HPC2 U3495 ( .a ({state_in_s1[72], state_in_s0[72]}), .b ({state_in_s1[264], state_in_s0[264]}), .c ({new_AGEMA_signal_2671, n3386}) ) ;
    xnor_HPC2 U3500 ( .a ({state_in_s1[75], state_in_s0[75]}), .b ({state_in_s1[267], state_in_s0[267]}), .c ({new_AGEMA_signal_2673, n3388}) ) ;
    xnor_HPC2 U3561 ( .a ({state_in_s1[76], state_in_s0[76]}), .b ({state_in_s1[268], state_in_s0[268]}), .c ({new_AGEMA_signal_2675, n3430}) ) ;
    xnor_HPC2 U3579 ( .a ({state_in_s1[115], state_in_s0[115]}), .b ({state_in_s1[307], state_in_s0[307]}), .c ({new_AGEMA_signal_2677, n3449}) ) ;
    xnor_HPC2 U3607 ( .a ({state_in_s1[100], state_in_s0[100]}), .b ({state_in_s1[292], state_in_s0[292]}), .c ({new_AGEMA_signal_2679, n3469}) ) ;
    xnor_HPC2 U3669 ( .a ({state_in_s1[101], state_in_s0[101]}), .b ({state_in_s1[293], state_in_s0[293]}), .c ({new_AGEMA_signal_2681, n3520}) ) ;
    xnor_HPC2 U3701 ( .a ({state_in_s1[110], state_in_s0[110]}), .b ({state_in_s1[302], state_in_s0[302]}), .c ({new_AGEMA_signal_2683, n3547}) ) ;
    xnor_HPC2 U3771 ( .a ({state_in_s1[81], state_in_s0[81]}), .b ({state_in_s1[273], state_in_s0[273]}), .c ({new_AGEMA_signal_2685, n3610}) ) ;
    xnor_HPC2 U3864 ( .a ({state_in_s1[84], state_in_s0[84]}), .b ({state_in_s1[276], state_in_s0[276]}), .c ({new_AGEMA_signal_2687, n3699}) ) ;
    xnor_HPC2 U3949 ( .a ({state_in_s1[85], state_in_s0[85]}), .b ({state_in_s1[277], state_in_s0[277]}), .c ({new_AGEMA_signal_2689, n3793}) ) ;
    xor_HPC2 U4057 ( .a ({state_in_s1[177], state_in_s0[177]}), .b ({state_in_s1[113], state_in_s0[113]}), .c ({new_AGEMA_signal_2692, n3291}) ) ;
    xor_HPC2 U4058 ( .a ({state_in_s1[171], state_in_s0[171]}), .b ({state_in_s1[107], state_in_s0[107]}), .c ({new_AGEMA_signal_2695, n3280}) ) ;
    xor_HPC2 U4059 ( .a ({state_in_s1[98], state_in_s0[98]}), .b ({state_in_s1[162], state_in_s0[162]}), .c ({new_AGEMA_signal_2698, n3273}) ) ;
    xor_HPC2 U4071 ( .a ({state_in_s1[172], state_in_s0[172]}), .b ({state_in_s1[108], state_in_s0[108]}), .c ({new_AGEMA_signal_2701, n3279}) ) ;
    xor_HPC2 U4072 ( .a ({state_in_s1[178], state_in_s0[178]}), .b ({state_in_s1[114], state_in_s0[114]}), .c ({new_AGEMA_signal_2704, n3290}) ) ;
    xor_HPC2 U4073 ( .a ({state_in_s1[99], state_in_s0[99]}), .b ({state_in_s1[163], state_in_s0[163]}), .c ({new_AGEMA_signal_2707, n3272}) ) ;
    xor_HPC2 U4085 ( .a ({state_in_s1[115], state_in_s0[115]}), .b ({state_in_s1[179], state_in_s0[179]}), .c ({new_AGEMA_signal_2709, n3289}) ) ;
    xor_HPC2 U4086 ( .a ({state_in_s1[109], state_in_s0[109]}), .b ({state_in_s1[173], state_in_s0[173]}), .c ({new_AGEMA_signal_2712, n3278}) ) ;
    xor_HPC2 U4087 ( .a ({state_in_s1[100], state_in_s0[100]}), .b ({state_in_s1[164], state_in_s0[164]}), .c ({new_AGEMA_signal_2714, n3271}) ) ;
    xor_HPC2 U4099 ( .a ({state_in_s1[180], state_in_s0[180]}), .b ({state_in_s1[116], state_in_s0[116]}), .c ({new_AGEMA_signal_2717, n3288}) ) ;
    xor_HPC2 U4100 ( .a ({state_in_s1[110], state_in_s0[110]}), .b ({state_in_s1[174], state_in_s0[174]}), .c ({new_AGEMA_signal_2719, n3277}) ) ;
    xor_HPC2 U4101 ( .a ({state_in_s1[101], state_in_s0[101]}), .b ({state_in_s1[165], state_in_s0[165]}), .c ({new_AGEMA_signal_2721, n3270}) ) ;
    xor_HPC2 U4113 ( .a ({state_in_s1[175], state_in_s0[175]}), .b ({state_in_s1[111], state_in_s0[111]}), .c ({new_AGEMA_signal_2724, n3276}) ) ;
    xor_HPC2 U4114 ( .a ({state_in_s1[181], state_in_s0[181]}), .b ({state_in_s1[117], state_in_s0[117]}), .c ({new_AGEMA_signal_2727, n3286}) ) ;
    xor_HPC2 U4115 ( .a ({state_in_s1[102], state_in_s0[102]}), .b ({state_in_s1[166], state_in_s0[166]}), .c ({new_AGEMA_signal_2730, n3269}) ) ;
    xor_HPC2 U4127 ( .a ({state_in_s1[182], state_in_s0[182]}), .b ({state_in_s1[118], state_in_s0[118]}), .c ({new_AGEMA_signal_2733, n3285}) ) ;
    xor_HPC2 U4128 ( .a ({state_in_s1[160], state_in_s0[160]}), .b ({state_in_s1[96], state_in_s0[96]}), .c ({new_AGEMA_signal_2736, n3275}) ) ;
    xor_HPC2 U4129 ( .a ({state_in_s1[103], state_in_s0[103]}), .b ({state_in_s1[167], state_in_s0[167]}), .c ({new_AGEMA_signal_2739, n3268}) ) ;
    xor_HPC2 U4141 ( .a ({state_in_s1[119], state_in_s0[119]}), .b ({state_in_s1[183], state_in_s0[183]}), .c ({new_AGEMA_signal_2742, n3284}) ) ;
    xor_HPC2 U4142 ( .a ({state_in_s1[97], state_in_s0[97]}), .b ({state_in_s1[161], state_in_s0[161]}), .c ({new_AGEMA_signal_2744, n3274}) ) ;
    xor_HPC2 U4143 ( .a ({state_in_s1[88], state_in_s0[88]}), .b ({state_in_s1[152], state_in_s0[152]}), .c ({new_AGEMA_signal_2747, n3267}) ) ;
    xor_HPC2 U4155 ( .a ({state_in_s1[168], state_in_s0[168]}), .b ({state_in_s1[104], state_in_s0[104]}), .c ({new_AGEMA_signal_2750, n3283}) ) ;
    xor_HPC2 U4156 ( .a ({state_in_s1[89], state_in_s0[89]}), .b ({state_in_s1[153], state_in_s0[153]}), .c ({new_AGEMA_signal_2753, n3266}) ) ;
    xor_HPC2 U4165 ( .a ({state_in_s1[169], state_in_s0[169]}), .b ({state_in_s1[105], state_in_s0[105]}), .c ({new_AGEMA_signal_2755, n3282}) ) ;
    xor_HPC2 U4166 ( .a ({state_in_s1[90], state_in_s0[90]}), .b ({state_in_s1[154], state_in_s0[154]}), .c ({new_AGEMA_signal_2758, n3265}) ) ;
    xor_HPC2 U4175 ( .a ({state_in_s1[106], state_in_s0[106]}), .b ({state_in_s1[170], state_in_s0[170]}), .c ({new_AGEMA_signal_2760, n3281}) ) ;
    xor_HPC2 U4176 ( .a ({state_in_s1[91], state_in_s0[91]}), .b ({state_in_s1[155], state_in_s0[155]}), .c ({new_AGEMA_signal_2763, n3264}) ) ;
    xor_HPC2 U4185 ( .a ({state_in_s1[92], state_in_s0[92]}), .b ({state_in_s1[156], state_in_s0[156]}), .c ({new_AGEMA_signal_2766, n3263}) ) ;
    xor_HPC2 U4191 ( .a ({state_in_s1[93], state_in_s0[93]}), .b ({state_in_s1[157], state_in_s0[157]}), .c ({new_AGEMA_signal_2769, n3262}) ) ;
    xor_HPC2 U4197 ( .a ({state_in_s1[94], state_in_s0[94]}), .b ({state_in_s1[158], state_in_s0[158]}), .c ({new_AGEMA_signal_2772, n3261}) ) ;
    xor_HPC2 U4203 ( .a ({state_in_s1[95], state_in_s0[95]}), .b ({state_in_s1[159], state_in_s0[159]}), .c ({new_AGEMA_signal_2775, n3260}) ) ;
    xor_HPC2 U4209 ( .a ({state_in_s1[80], state_in_s0[80]}), .b ({state_in_s1[144], state_in_s0[144]}), .c ({new_AGEMA_signal_2778, n3259}) ) ;
    xor_HPC2 U4215 ( .a ({state_in_s1[81], state_in_s0[81]}), .b ({state_in_s1[145], state_in_s0[145]}), .c ({new_AGEMA_signal_2780, n3258}) ) ;
    xor_HPC2 U4221 ( .a ({state_in_s1[82], state_in_s0[82]}), .b ({state_in_s1[146], state_in_s0[146]}), .c ({new_AGEMA_signal_2783, n3257}) ) ;
    xor_HPC2 U4227 ( .a ({state_in_s1[83], state_in_s0[83]}), .b ({state_in_s1[147], state_in_s0[147]}), .c ({new_AGEMA_signal_2786, n3256}) ) ;
    xor_HPC2 U4233 ( .a ({state_in_s1[84], state_in_s0[84]}), .b ({state_in_s1[148], state_in_s0[148]}), .c ({new_AGEMA_signal_2788, n3255}) ) ;
    xor_HPC2 U4239 ( .a ({state_in_s1[85], state_in_s0[85]}), .b ({state_in_s1[149], state_in_s0[149]}), .c ({new_AGEMA_signal_2790, n3254}) ) ;
    xor_HPC2 U4245 ( .a ({state_in_s1[86], state_in_s0[86]}), .b ({state_in_s1[150], state_in_s0[150]}), .c ({new_AGEMA_signal_2793, n3253}) ) ;
    xor_HPC2 U4251 ( .a ({state_in_s1[87], state_in_s0[87]}), .b ({state_in_s1[151], state_in_s0[151]}), .c ({new_AGEMA_signal_2795, n3252}) ) ;
    xor_HPC2 U4257 ( .a ({state_in_s1[72], state_in_s0[72]}), .b ({state_in_s1[136], state_in_s0[136]}), .c ({new_AGEMA_signal_2797, n3251}) ) ;
    xor_HPC2 U4263 ( .a ({state_in_s1[137], state_in_s0[137]}), .b ({state_in_s1[73], state_in_s0[73]}), .c ({new_AGEMA_signal_2800, n3250}) ) ;
    xor_HPC2 U4269 ( .a ({state_in_s1[138], state_in_s0[138]}), .b ({state_in_s1[74], state_in_s0[74]}), .c ({new_AGEMA_signal_2803, n3249}) ) ;
    xor_HPC2 U4275 ( .a ({state_in_s1[75], state_in_s0[75]}), .b ({state_in_s1[139], state_in_s0[139]}), .c ({new_AGEMA_signal_2805, n3248}) ) ;
    xor_HPC2 U4281 ( .a ({state_in_s1[76], state_in_s0[76]}), .b ({state_in_s1[140], state_in_s0[140]}), .c ({new_AGEMA_signal_2807, n3247}) ) ;
    xor_HPC2 U4287 ( .a ({state_in_s1[141], state_in_s0[141]}), .b ({state_in_s1[77], state_in_s0[77]}), .c ({new_AGEMA_signal_2810, n3246}) ) ;
    xor_HPC2 U4293 ( .a ({state_in_s1[142], state_in_s0[142]}), .b ({state_in_s1[78], state_in_s0[78]}), .c ({new_AGEMA_signal_2813, n3245}) ) ;
    xor_HPC2 U4299 ( .a ({state_in_s1[79], state_in_s0[79]}), .b ({state_in_s1[143], state_in_s0[143]}), .c ({new_AGEMA_signal_2816, n3244}) ) ;
    xor_HPC2 U4305 ( .a ({state_in_s1[128], state_in_s0[128]}), .b ({state_in_s1[64], state_in_s0[64]}), .c ({new_AGEMA_signal_2819, n3243}) ) ;
    xor_HPC2 U4311 ( .a ({state_in_s1[129], state_in_s0[129]}), .b ({state_in_s1[65], state_in_s0[65]}), .c ({new_AGEMA_signal_2821, n3242}) ) ;
    xor_HPC2 U4317 ( .a ({state_in_s1[66], state_in_s0[66]}), .b ({state_in_s1[130], state_in_s0[130]}), .c ({new_AGEMA_signal_2823, n3241}) ) ;
    xor_HPC2 U4323 ( .a ({state_in_s1[131], state_in_s0[131]}), .b ({state_in_s1[67], state_in_s0[67]}), .c ({new_AGEMA_signal_2825, n3240}) ) ;
    xor_HPC2 U4329 ( .a ({state_in_s1[132], state_in_s0[132]}), .b ({state_in_s1[68], state_in_s0[68]}), .c ({new_AGEMA_signal_2828, n3238}) ) ;
    xor_HPC2 U4335 ( .a ({state_in_s1[184], state_in_s0[184]}), .b ({state_in_s1[120], state_in_s0[120]}), .c ({new_AGEMA_signal_2831, n4041}) ) ;
    INV_X1 U4344 ( .A (rcon[0]), .ZN (n4068) ) ;
    xnor_HPC2 U4345 ( .a ({new_AGEMA_signal_2831, n4041}), .b ({1'b0, n4068}), .c ({new_AGEMA_signal_2989, y2[0]}) ) ;
    xor_HPC2 U4346 ( .a ({state_in_s1[176], state_in_s0[176]}), .b ({state_in_s1[112], state_in_s0[112]}), .c ({new_AGEMA_signal_2834, n3237}) ) ;
    xor_HPC2 U4352 ( .a ({state_in_s1[133], state_in_s0[133]}), .b ({state_in_s1[69], state_in_s0[69]}), .c ({new_AGEMA_signal_2837, n3236}) ) ;
    xor_HPC2 U4358 ( .a ({state_in_s1[134], state_in_s0[134]}), .b ({state_in_s1[70], state_in_s0[70]}), .c ({new_AGEMA_signal_2840, n3235}) ) ;
    xor_HPC2 U4366 ( .a ({state_in_s1[188], state_in_s0[188]}), .b ({state_in_s1[124], state_in_s0[124]}), .c ({new_AGEMA_signal_2843, n4208}) ) ;
    xnor_HPC2 U4367 ( .a ({1'b0, rcon[0]}), .b ({new_AGEMA_signal_2843, n4208}), .c ({new_AGEMA_signal_2990, n3232}) ) ;
    xor_HPC2 U4368 ( .a ({state_in_s1[135], state_in_s0[135]}), .b ({state_in_s1[71], state_in_s0[71]}), .c ({new_AGEMA_signal_2846, n3234}) ) ;
    INV_X1 U4379 ( .A (rcon[1]), .ZN (n4067) ) ;
    XNOR2_X1 U4380 ( .A (rcon[0]), .B (n4067), .ZN (n4206) ) ;
    xor_HPC2 U4381 ( .a ({state_in_s1[185], state_in_s0[185]}), .b ({state_in_s1[121], state_in_s0[121]}), .c ({new_AGEMA_signal_2849, n4066}) ) ;
    xor_HPC2 U4392 ( .a ({1'b0, n4206}), .b ({new_AGEMA_signal_2849, n4066}), .c ({new_AGEMA_signal_3513, y2[1]}) ) ;
    xnor_HPC2 U4393 ( .a ({state_in_s1[186], state_in_s0[186]}), .b ({state_in_s1[122], state_in_s0[122]}), .c ({new_AGEMA_signal_2852, n4069}) ) ;
    NAND2_X1 U4394 ( .A1 (n4068), .A2 (n4067), .ZN (n4079) ) ;
    XNOR2_X1 U4395 ( .A (rcon[2]), .B (n4079), .ZN (n4087) ) ;
    xnor_HPC2 U4396 ( .a ({new_AGEMA_signal_2852, n4069}), .b ({1'b0, n4087}), .c ({new_AGEMA_signal_3824, n3287}) ) ;
    NAND2_X1 U4406 ( .A1 (rcon[2]), .A2 (n4079), .ZN (n4080) ) ;
    XNOR2_X1 U4407 ( .A (rcon[3]), .B (n4080), .ZN (n4084) ) ;
    xor_HPC2 U4408 ( .a ({1'b0, n4084}), .b ({state_in_s1[187], state_in_s0[187]}), .c ({new_AGEMA_signal_4140, n4081}) ) ;
    xnor_HPC2 U4409 ( .a ({state_in_s1[123], state_in_s0[123]}), .b ({new_AGEMA_signal_4140, n4081}), .c ({new_AGEMA_signal_4432, n3233}) ) ;
    xnor_HPC2 U4415 ( .a ({1'b0, n4084}), .b ({state_in_s1[191], state_in_s0[191]}), .c ({new_AGEMA_signal_4142, n4085}) ) ;
    xnor_HPC2 U4416 ( .a ({new_AGEMA_signal_4142, n4085}), .b ({state_in_s1[127], state_in_s0[127]}), .c ({new_AGEMA_signal_4433, n3239}) ) ;
    xor_HPC2 U4417 ( .a ({state_in_s1[190], state_in_s0[190]}), .b ({state_in_s1[126], state_in_s0[126]}), .c ({new_AGEMA_signal_2855, n4086}) ) ;
    xnor_HPC2 U4418 ( .a ({1'b0, n4087}), .b ({new_AGEMA_signal_2855, n4086}), .c ({new_AGEMA_signal_3826, n3230}) ) ;
    xnor_HPC2 U4432 ( .a ({state_in_s1[125], state_in_s0[125]}), .b ({state_in_s1[189], state_in_s0[189]}), .c ({new_AGEMA_signal_2858, n4103}) ) ;
    xor_HPC2 U4439 ( .a ({1'b0, n4206}), .b ({new_AGEMA_signal_2858, n4103}), .c ({new_AGEMA_signal_3515, n3231}) ) ;
    not_masked SboxInst_U447 ( .a ({new_AGEMA_signal_2655, y0[0]}), .b ({new_AGEMA_signal_3047, SboxInst_n320}) ) ;
    not_masked SboxInst_U445 ( .a ({new_AGEMA_signal_2653, y0[10]}), .b ({new_AGEMA_signal_3048, SboxInst_n319}) ) ;
    not_masked SboxInst_U443 ( .a ({new_AGEMA_signal_2651, y0[11]}), .b ({new_AGEMA_signal_3049, SboxInst_n318}) ) ;
    not_masked SboxInst_U441 ( .a ({new_AGEMA_signal_2649, y0[12]}), .b ({new_AGEMA_signal_3050, SboxInst_n317}) ) ;
    not_masked SboxInst_U439 ( .a ({new_AGEMA_signal_2647, y0[13]}), .b ({new_AGEMA_signal_3051, SboxInst_n316}) ) ;
    not_masked SboxInst_U437 ( .a ({new_AGEMA_signal_2645, y0[14]}), .b ({new_AGEMA_signal_3052, SboxInst_n315}) ) ;
    not_masked SboxInst_U435 ( .a ({new_AGEMA_signal_2643, y0[15]}), .b ({new_AGEMA_signal_3053, SboxInst_n314}) ) ;
    not_masked SboxInst_U433 ( .a ({new_AGEMA_signal_2641, y0[16]}), .b ({new_AGEMA_signal_3054, SboxInst_n313}) ) ;
    not_masked SboxInst_U431 ( .a ({new_AGEMA_signal_2639, y0[17]}), .b ({new_AGEMA_signal_3055, SboxInst_n312}) ) ;
    not_masked SboxInst_U429 ( .a ({new_AGEMA_signal_2637, y0[18]}), .b ({new_AGEMA_signal_3056, SboxInst_n311}) ) ;
    not_masked SboxInst_U427 ( .a ({new_AGEMA_signal_2635, y0[19]}), .b ({new_AGEMA_signal_3057, SboxInst_n310}) ) ;
    not_masked SboxInst_U425 ( .a ({new_AGEMA_signal_2633, y0[1]}), .b ({new_AGEMA_signal_3058, SboxInst_n309}) ) ;
    not_masked SboxInst_U423 ( .a ({new_AGEMA_signal_2631, y0[20]}), .b ({new_AGEMA_signal_3059, SboxInst_n308}) ) ;
    not_masked SboxInst_U421 ( .a ({new_AGEMA_signal_2629, y0[21]}), .b ({new_AGEMA_signal_3060, SboxInst_n307}) ) ;
    not_masked SboxInst_U419 ( .a ({new_AGEMA_signal_2627, y0[22]}), .b ({new_AGEMA_signal_3061, SboxInst_n306}) ) ;
    not_masked SboxInst_U417 ( .a ({new_AGEMA_signal_2625, y0[23]}), .b ({new_AGEMA_signal_3062, SboxInst_n305}) ) ;
    not_masked SboxInst_U415 ( .a ({new_AGEMA_signal_2623, y0[24]}), .b ({new_AGEMA_signal_3063, SboxInst_n304}) ) ;
    not_masked SboxInst_U413 ( .a ({new_AGEMA_signal_2621, y0[25]}), .b ({new_AGEMA_signal_3064, SboxInst_n303}) ) ;
    not_masked SboxInst_U411 ( .a ({new_AGEMA_signal_2619, y0[26]}), .b ({new_AGEMA_signal_3065, SboxInst_n302}) ) ;
    not_masked SboxInst_U409 ( .a ({new_AGEMA_signal_2617, y0[27]}), .b ({new_AGEMA_signal_3066, SboxInst_n301}) ) ;
    not_masked SboxInst_U407 ( .a ({new_AGEMA_signal_2615, y0[28]}), .b ({new_AGEMA_signal_3067, SboxInst_n300}) ) ;
    not_masked SboxInst_U405 ( .a ({new_AGEMA_signal_2613, y0[29]}), .b ({new_AGEMA_signal_3068, SboxInst_n299}) ) ;
    not_masked SboxInst_U403 ( .a ({new_AGEMA_signal_2611, y0[2]}), .b ({new_AGEMA_signal_3069, SboxInst_n298}) ) ;
    not_masked SboxInst_U401 ( .a ({new_AGEMA_signal_2609, y0[30]}), .b ({new_AGEMA_signal_3070, SboxInst_n297}) ) ;
    not_masked SboxInst_U399 ( .a ({new_AGEMA_signal_2607, y0[31]}), .b ({new_AGEMA_signal_3071, SboxInst_n296}) ) ;
    not_masked SboxInst_U397 ( .a ({new_AGEMA_signal_2605, y0[32]}), .b ({new_AGEMA_signal_3072, SboxInst_n295}) ) ;
    not_masked SboxInst_U395 ( .a ({new_AGEMA_signal_2603, y0[33]}), .b ({new_AGEMA_signal_3073, SboxInst_n294}) ) ;
    not_masked SboxInst_U393 ( .a ({new_AGEMA_signal_2601, y0[34]}), .b ({new_AGEMA_signal_3074, SboxInst_n293}) ) ;
    not_masked SboxInst_U391 ( .a ({new_AGEMA_signal_2599, y0[35]}), .b ({new_AGEMA_signal_3075, SboxInst_n292}) ) ;
    not_masked SboxInst_U389 ( .a ({new_AGEMA_signal_2597, y0[36]}), .b ({new_AGEMA_signal_3076, SboxInst_n291}) ) ;
    not_masked SboxInst_U387 ( .a ({new_AGEMA_signal_2595, y0[37]}), .b ({new_AGEMA_signal_3077, SboxInst_n290}) ) ;
    not_masked SboxInst_U385 ( .a ({new_AGEMA_signal_2593, y0[38]}), .b ({new_AGEMA_signal_3078, SboxInst_n289}) ) ;
    not_masked SboxInst_U383 ( .a ({new_AGEMA_signal_2591, y0[39]}), .b ({new_AGEMA_signal_3079, SboxInst_n288}) ) ;
    not_masked SboxInst_U381 ( .a ({new_AGEMA_signal_2589, y0[3]}), .b ({new_AGEMA_signal_3080, SboxInst_n287}) ) ;
    not_masked SboxInst_U379 ( .a ({new_AGEMA_signal_2587, y0[40]}), .b ({new_AGEMA_signal_3081, SboxInst_n286}) ) ;
    not_masked SboxInst_U377 ( .a ({new_AGEMA_signal_2585, y0[41]}), .b ({new_AGEMA_signal_3082, SboxInst_n285}) ) ;
    not_masked SboxInst_U375 ( .a ({new_AGEMA_signal_2583, y0[42]}), .b ({new_AGEMA_signal_3083, SboxInst_n284}) ) ;
    not_masked SboxInst_U373 ( .a ({new_AGEMA_signal_2581, y0[43]}), .b ({new_AGEMA_signal_3084, SboxInst_n283}) ) ;
    not_masked SboxInst_U371 ( .a ({new_AGEMA_signal_2579, y0[44]}), .b ({new_AGEMA_signal_3085, SboxInst_n282}) ) ;
    not_masked SboxInst_U369 ( .a ({new_AGEMA_signal_2577, y0[45]}), .b ({new_AGEMA_signal_3086, SboxInst_n281}) ) ;
    not_masked SboxInst_U367 ( .a ({new_AGEMA_signal_2575, y0[46]}), .b ({new_AGEMA_signal_3087, SboxInst_n280}) ) ;
    not_masked SboxInst_U365 ( .a ({new_AGEMA_signal_2573, y0[47]}), .b ({new_AGEMA_signal_3088, SboxInst_n279}) ) ;
    not_masked SboxInst_U363 ( .a ({new_AGEMA_signal_2571, y0[48]}), .b ({new_AGEMA_signal_3089, SboxInst_n278}) ) ;
    not_masked SboxInst_U361 ( .a ({new_AGEMA_signal_2569, y0[49]}), .b ({new_AGEMA_signal_3090, SboxInst_n277}) ) ;
    not_masked SboxInst_U359 ( .a ({new_AGEMA_signal_2567, y0[4]}), .b ({new_AGEMA_signal_3091, SboxInst_n276}) ) ;
    not_masked SboxInst_U357 ( .a ({new_AGEMA_signal_2565, y0[50]}), .b ({new_AGEMA_signal_3092, SboxInst_n275}) ) ;
    not_masked SboxInst_U355 ( .a ({new_AGEMA_signal_2563, y0[51]}), .b ({new_AGEMA_signal_3093, SboxInst_n274}) ) ;
    not_masked SboxInst_U353 ( .a ({new_AGEMA_signal_2561, y0[52]}), .b ({new_AGEMA_signal_3094, SboxInst_n273}) ) ;
    not_masked SboxInst_U351 ( .a ({new_AGEMA_signal_2559, y0[53]}), .b ({new_AGEMA_signal_3095, SboxInst_n272}) ) ;
    not_masked SboxInst_U349 ( .a ({new_AGEMA_signal_2557, y0[54]}), .b ({new_AGEMA_signal_3096, SboxInst_n271}) ) ;
    not_masked SboxInst_U347 ( .a ({new_AGEMA_signal_2555, y0[55]}), .b ({new_AGEMA_signal_3097, SboxInst_n270}) ) ;
    not_masked SboxInst_U345 ( .a ({new_AGEMA_signal_2553, y0[56]}), .b ({new_AGEMA_signal_3098, SboxInst_n269}) ) ;
    not_masked SboxInst_U343 ( .a ({new_AGEMA_signal_2551, y0[57]}), .b ({new_AGEMA_signal_3099, SboxInst_n268}) ) ;
    not_masked SboxInst_U341 ( .a ({new_AGEMA_signal_2549, y0[58]}), .b ({new_AGEMA_signal_3100, SboxInst_n267}) ) ;
    not_masked SboxInst_U339 ( .a ({new_AGEMA_signal_2547, y0[59]}), .b ({new_AGEMA_signal_3101, SboxInst_n266}) ) ;
    not_masked SboxInst_U337 ( .a ({new_AGEMA_signal_2545, y0[5]}), .b ({new_AGEMA_signal_3102, SboxInst_n265}) ) ;
    not_masked SboxInst_U335 ( .a ({new_AGEMA_signal_2543, y0[60]}), .b ({new_AGEMA_signal_3103, SboxInst_n264}) ) ;
    not_masked SboxInst_U333 ( .a ({new_AGEMA_signal_2541, y0[61]}), .b ({new_AGEMA_signal_3104, SboxInst_n263}) ) ;
    not_masked SboxInst_U331 ( .a ({new_AGEMA_signal_2539, y0[62]}), .b ({new_AGEMA_signal_3105, SboxInst_n262}) ) ;
    not_masked SboxInst_U329 ( .a ({new_AGEMA_signal_2537, y0[63]}), .b ({new_AGEMA_signal_3106, SboxInst_n261}) ) ;
    not_masked SboxInst_U327 ( .a ({new_AGEMA_signal_2535, y0[6]}), .b ({new_AGEMA_signal_3107, SboxInst_n260}) ) ;
    not_masked SboxInst_U325 ( .a ({new_AGEMA_signal_2533, y0[7]}), .b ({new_AGEMA_signal_3108, SboxInst_n259}) ) ;
    not_masked SboxInst_U323 ( .a ({new_AGEMA_signal_2531, y0[8]}), .b ({new_AGEMA_signal_3109, SboxInst_n258}) ) ;
    not_masked SboxInst_U321 ( .a ({new_AGEMA_signal_2529, y0[9]}), .b ({new_AGEMA_signal_3110, SboxInst_n257}) ) ;
    not_masked SboxInst_U255 ( .a ({state_in_s1[213], state_in_s0[213]}), .b ({new_AGEMA_signal_2859, SboxInst_n345}) ) ;
    not_masked SboxInst_U253 ( .a ({state_in_s1[223], state_in_s0[223]}), .b ({new_AGEMA_signal_2860, SboxInst_n352}) ) ;
    not_masked SboxInst_U251 ( .a ({state_in_s1[208], state_in_s0[208]}), .b ({new_AGEMA_signal_2861, SboxInst_n350}) ) ;
    not_masked SboxInst_U249 ( .a ({state_in_s1[212], state_in_s0[212]}), .b ({new_AGEMA_signal_2862, SboxInst_n346}) ) ;
    not_masked SboxInst_U247 ( .a ({state_in_s1[222], state_in_s0[222]}), .b ({new_AGEMA_signal_2863, SboxInst_n353}) ) ;
    not_masked SboxInst_U245 ( .a ({state_in_s1[211], state_in_s0[211]}), .b ({new_AGEMA_signal_2864, SboxInst_n347}) ) ;
    not_masked SboxInst_U243 ( .a ({state_in_s1[221], state_in_s0[221]}), .b ({new_AGEMA_signal_2865, SboxInst_n354}) ) ;
    not_masked SboxInst_U241 ( .a ({state_in_s1[210], state_in_s0[210]}), .b ({new_AGEMA_signal_2866, SboxInst_n348}) ) ;
    not_masked SboxInst_U239 ( .a ({state_in_s1[220], state_in_s0[220]}), .b ({new_AGEMA_signal_2867, SboxInst_n355}) ) ;
    not_masked SboxInst_U237 ( .a ({state_in_s1[209], state_in_s0[209]}), .b ({new_AGEMA_signal_2868, SboxInst_n349}) ) ;
    not_masked SboxInst_U235 ( .a ({state_in_s1[219], state_in_s0[219]}), .b ({new_AGEMA_signal_2869, SboxInst_n356}) ) ;
    not_masked SboxInst_U233 ( .a ({state_in_s1[218], state_in_s0[218]}), .b ({new_AGEMA_signal_2870, SboxInst_n357}) ) ;
    not_masked SboxInst_U231 ( .a ({state_in_s1[217], state_in_s0[217]}), .b ({new_AGEMA_signal_2871, SboxInst_n358}) ) ;
    not_masked SboxInst_U229 ( .a ({state_in_s1[216], state_in_s0[216]}), .b ({new_AGEMA_signal_2872, SboxInst_n359}) ) ;
    not_masked SboxInst_U227 ( .a ({state_in_s1[200], state_in_s0[200]}), .b ({new_AGEMA_signal_2873, SboxInst_n342}) ) ;
    not_masked SboxInst_U225 ( .a ({state_in_s1[205], state_in_s0[205]}), .b ({new_AGEMA_signal_2874, SboxInst_n336}) ) ;
    not_masked SboxInst_U223 ( .a ({state_in_s1[215], state_in_s0[215]}), .b ({new_AGEMA_signal_2875, SboxInst_n343}) ) ;
    not_masked SboxInst_U221 ( .a ({state_in_s1[204], state_in_s0[204]}), .b ({new_AGEMA_signal_2876, SboxInst_n337}) ) ;
    not_masked SboxInst_U219 ( .a ({state_in_s1[214], state_in_s0[214]}), .b ({new_AGEMA_signal_2877, SboxInst_n344}) ) ;
    not_masked SboxInst_U217 ( .a ({state_in_s1[203], state_in_s0[203]}), .b ({new_AGEMA_signal_2878, SboxInst_n338}) ) ;
    not_masked SboxInst_U215 ( .a ({state_in_s1[202], state_in_s0[202]}), .b ({new_AGEMA_signal_2879, SboxInst_n339}) ) ;
    not_masked SboxInst_U213 ( .a ({state_in_s1[201], state_in_s0[201]}), .b ({new_AGEMA_signal_2880, SboxInst_n341}) ) ;
    not_masked SboxInst_U211 ( .a ({state_in_s1[207], state_in_s0[207]}), .b ({new_AGEMA_signal_2881, SboxInst_n334}) ) ;
    not_masked SboxInst_U209 ( .a ({state_in_s1[197], state_in_s0[197]}), .b ({new_AGEMA_signal_2882, SboxInst_n327}) ) ;
    not_masked SboxInst_U207 ( .a ({state_in_s1[192], state_in_s0[192]}), .b ({new_AGEMA_signal_2883, SboxInst_n333}) ) ;
    not_masked SboxInst_U205 ( .a ({state_in_s1[206], state_in_s0[206]}), .b ({new_AGEMA_signal_2884, SboxInst_n335}) ) ;
    not_masked SboxInst_U203 ( .a ({state_in_s1[196], state_in_s0[196]}), .b ({new_AGEMA_signal_2885, SboxInst_n328}) ) ;
    not_masked SboxInst_U201 ( .a ({state_in_s1[195], state_in_s0[195]}), .b ({new_AGEMA_signal_2886, SboxInst_n330}) ) ;
    not_masked SboxInst_U199 ( .a ({state_in_s1[194], state_in_s0[194]}), .b ({new_AGEMA_signal_2887, SboxInst_n331}) ) ;
    not_masked SboxInst_U197 ( .a ({state_in_s1[193], state_in_s0[193]}), .b ({new_AGEMA_signal_2888, SboxInst_n332}) ) ;
    not_masked SboxInst_U195 ( .a ({state_in_s1[199], state_in_s0[199]}), .b ({new_AGEMA_signal_2889, SboxInst_n325}) ) ;
    not_masked SboxInst_U193 ( .a ({state_in_s1[248], state_in_s0[248]}), .b ({new_AGEMA_signal_2890, SboxInst_n384}) ) ;
    not_masked SboxInst_U191 ( .a ({state_in_s1[253], state_in_s0[253]}), .b ({new_AGEMA_signal_2891, SboxInst_n329}) ) ;
    not_masked SboxInst_U189 ( .a ({state_in_s1[252], state_in_s0[252]}), .b ({new_AGEMA_signal_2892, SboxInst_n340}) ) ;
    not_masked SboxInst_U187 ( .a ({state_in_s1[198], state_in_s0[198]}), .b ({new_AGEMA_signal_2893, SboxInst_n326}) ) ;
    not_masked SboxInst_U185 ( .a ({state_in_s1[251], state_in_s0[251]}), .b ({new_AGEMA_signal_2894, SboxInst_n351}) ) ;
    not_masked SboxInst_U183 ( .a ({state_in_s1[250], state_in_s0[250]}), .b ({new_AGEMA_signal_2895, SboxInst_n362}) ) ;
    not_masked SboxInst_U181 ( .a ({state_in_s1[249], state_in_s0[249]}), .b ({new_AGEMA_signal_2896, SboxInst_n373}) ) ;
    not_masked SboxInst_U179 ( .a ({state_in_s1[86], state_in_s0[86]}), .b ({new_AGEMA_signal_2897, SboxInst_n216}) ) ;
    not_masked SboxInst_U177 ( .a ({state_in_s1[127], state_in_s0[127]}), .b ({new_AGEMA_signal_2899, SboxInst_n195}) ) ;
    not_masked SboxInst_U175 ( .a ({state_in_s1[124], state_in_s0[124]}), .b ({new_AGEMA_signal_2900, SboxInst_n212}) ) ;
    not_masked SboxInst_U173 ( .a ({state_in_s1[126], state_in_s0[126]}), .b ({new_AGEMA_signal_2901, SboxInst_n196}) ) ;
    not_masked SboxInst_U171 ( .a ({state_in_s1[85], state_in_s0[85]}), .b ({new_AGEMA_signal_2902, SboxInst_n217}) ) ;
    not_masked SboxInst_U169 ( .a ({state_in_s1[123], state_in_s0[123]}), .b ({new_AGEMA_signal_2904, SboxInst_n223}) ) ;
    not_masked SboxInst_U167 ( .a ({state_in_s1[84], state_in_s0[84]}), .b ({new_AGEMA_signal_2905, SboxInst_n218}) ) ;
    not_masked SboxInst_U165 ( .a ({state_in_s1[122], state_in_s0[122]}), .b ({new_AGEMA_signal_2906, SboxInst_n234}) ) ;
    not_masked SboxInst_U163 ( .a ({state_in_s1[125], state_in_s0[125]}), .b ({new_AGEMA_signal_2907, SboxInst_n201}) ) ;
    not_masked SboxInst_U161 ( .a ({state_in_s1[83], state_in_s0[83]}), .b ({new_AGEMA_signal_2908, SboxInst_n219}) ) ;
    not_masked SboxInst_U159 ( .a ({state_in_s1[121], state_in_s0[121]}), .b ({new_AGEMA_signal_2909, SboxInst_n245}) ) ;
    not_masked SboxInst_U157 ( .a ({state_in_s1[82], state_in_s0[82]}), .b ({new_AGEMA_signal_2910, SboxInst_n220}) ) ;
    not_masked SboxInst_U155 ( .a ({state_in_s1[120], state_in_s0[120]}), .b ({new_AGEMA_signal_2911, SboxInst_n256}) ) ;
    not_masked SboxInst_U153 ( .a ({state_in_s1[71], state_in_s0[71]}), .b ({new_AGEMA_signal_2912, SboxInst_n197}) ) ;
    not_masked SboxInst_U151 ( .a ({state_in_s1[81], state_in_s0[81]}), .b ({new_AGEMA_signal_2913, SboxInst_n221}) ) ;
    not_masked SboxInst_U149 ( .a ({state_in_s1[80], state_in_s0[80]}), .b ({new_AGEMA_signal_2914, SboxInst_n222}) ) ;
    not_masked SboxInst_U147 ( .a ({state_in_s1[70], state_in_s0[70]}), .b ({new_AGEMA_signal_2915, SboxInst_n198}) ) ;
    not_masked SboxInst_U145 ( .a ({state_in_s1[95], state_in_s0[95]}), .b ({new_AGEMA_signal_2916, SboxInst_n224}) ) ;
    not_masked SboxInst_U143 ( .a ({state_in_s1[69], state_in_s0[69]}), .b ({new_AGEMA_signal_2917, SboxInst_n199}) ) ;
    not_masked SboxInst_U141 ( .a ({state_in_s1[119], state_in_s0[119]}), .b ({new_AGEMA_signal_2918, SboxInst_n250}) ) ;
    not_masked SboxInst_U139 ( .a ({state_in_s1[116], state_in_s0[116]}), .b ({new_AGEMA_signal_2919, SboxInst_n253}) ) ;
    not_masked SboxInst_U137 ( .a ({state_in_s1[78], state_in_s0[78]}), .b ({new_AGEMA_signal_2920, SboxInst_n207}) ) ;
    not_masked SboxInst_U135 ( .a ({state_in_s1[115], state_in_s0[115]}), .b ({new_AGEMA_signal_2921, SboxInst_n254}) ) ;
    not_masked SboxInst_U133 ( .a ({state_in_s1[118], state_in_s0[118]}), .b ({new_AGEMA_signal_2922, SboxInst_n251}) ) ;
    not_masked SboxInst_U131 ( .a ({state_in_s1[77], state_in_s0[77]}), .b ({new_AGEMA_signal_2923, SboxInst_n208}) ) ;
    not_masked SboxInst_U129 ( .a ({state_in_s1[114], state_in_s0[114]}), .b ({new_AGEMA_signal_2924, SboxInst_n255}) ) ;
    not_masked SboxInst_U127 ( .a ({state_in_s1[117], state_in_s0[117]}), .b ({new_AGEMA_signal_2925, SboxInst_n252}) ) ;
    not_masked SboxInst_U125 ( .a ({state_in_s1[76], state_in_s0[76]}), .b ({new_AGEMA_signal_2926, SboxInst_n209}) ) ;
    not_masked SboxInst_U123 ( .a ({state_in_s1[113], state_in_s0[113]}), .b ({new_AGEMA_signal_2927, SboxInst_n193}) ) ;
    not_masked SboxInst_U121 ( .a ({state_in_s1[75], state_in_s0[75]}), .b ({new_AGEMA_signal_2928, SboxInst_n210}) ) ;
    not_masked SboxInst_U119 ( .a ({state_in_s1[112], state_in_s0[112]}), .b ({new_AGEMA_signal_2929, SboxInst_n194}) ) ;
    not_masked SboxInst_U117 ( .a ({state_in_s1[74], state_in_s0[74]}), .b ({new_AGEMA_signal_2930, SboxInst_n211}) ) ;
    not_masked SboxInst_U115 ( .a ({state_in_s1[73], state_in_s0[73]}), .b ({new_AGEMA_signal_2931, SboxInst_n213}) ) ;
    not_masked SboxInst_U113 ( .a ({state_in_s1[72], state_in_s0[72]}), .b ({new_AGEMA_signal_2932, SboxInst_n214}) ) ;
    not_masked SboxInst_U111 ( .a ({state_in_s1[87], state_in_s0[87]}), .b ({new_AGEMA_signal_2933, SboxInst_n215}) ) ;
    not_masked SboxInst_U109 ( .a ({state_in_s1[108], state_in_s0[108]}), .b ({new_AGEMA_signal_2934, SboxInst_n244}) ) ;
    not_masked SboxInst_U107 ( .a ({state_in_s1[111], state_in_s0[111]}), .b ({new_AGEMA_signal_2935, SboxInst_n241}) ) ;
    not_masked SboxInst_U105 ( .a ({state_in_s1[107], state_in_s0[107]}), .b ({new_AGEMA_signal_2936, SboxInst_n246}) ) ;
    not_masked SboxInst_U103 ( .a ({state_in_s1[110], state_in_s0[110]}), .b ({new_AGEMA_signal_2937, SboxInst_n242}) ) ;
    not_masked SboxInst_U101 ( .a ({state_in_s1[68], state_in_s0[68]}), .b ({new_AGEMA_signal_2938, SboxInst_n200}) ) ;
    not_masked SboxInst_U99 ( .a ({state_in_s1[109], state_in_s0[109]}), .b ({new_AGEMA_signal_2939, SboxInst_n243}) ) ;
    not_masked SboxInst_U97 ( .a ({state_in_s1[106], state_in_s0[106]}), .b ({new_AGEMA_signal_2940, SboxInst_n247}) ) ;
    not_masked SboxInst_U95 ( .a ({state_in_s1[67], state_in_s0[67]}), .b ({new_AGEMA_signal_2941, SboxInst_n202}) ) ;
    not_masked SboxInst_U93 ( .a ({state_in_s1[105], state_in_s0[105]}), .b ({new_AGEMA_signal_2942, SboxInst_n248}) ) ;
    not_masked SboxInst_U91 ( .a ({state_in_s1[66], state_in_s0[66]}), .b ({new_AGEMA_signal_2943, SboxInst_n203}) ) ;
    not_masked SboxInst_U89 ( .a ({state_in_s1[104], state_in_s0[104]}), .b ({new_AGEMA_signal_2944, SboxInst_n249}) ) ;
    not_masked SboxInst_U87 ( .a ({state_in_s1[65], state_in_s0[65]}), .b ({new_AGEMA_signal_2945, SboxInst_n204}) ) ;
    not_masked SboxInst_U85 ( .a ({state_in_s1[64], state_in_s0[64]}), .b ({new_AGEMA_signal_2946, SboxInst_n205}) ) ;
    not_masked SboxInst_U83 ( .a ({state_in_s1[79], state_in_s0[79]}), .b ({new_AGEMA_signal_2947, SboxInst_n206}) ) ;
    not_masked SboxInst_U81 ( .a ({state_in_s1[103], state_in_s0[103]}), .b ({new_AGEMA_signal_2948, SboxInst_n232}) ) ;
    not_masked SboxInst_U79 ( .a ({state_in_s1[100], state_in_s0[100]}), .b ({new_AGEMA_signal_2949, SboxInst_n236}) ) ;
    not_masked SboxInst_U77 ( .a ({state_in_s1[102], state_in_s0[102]}), .b ({new_AGEMA_signal_2950, SboxInst_n233}) ) ;
    not_masked SboxInst_U75 ( .a ({state_in_s1[99], state_in_s0[99]}), .b ({new_AGEMA_signal_2951, SboxInst_n237}) ) ;
    not_masked SboxInst_U73 ( .a ({state_in_s1[98], state_in_s0[98]}), .b ({new_AGEMA_signal_2952, SboxInst_n238}) ) ;
    not_masked SboxInst_U71 ( .a ({state_in_s1[101], state_in_s0[101]}), .b ({new_AGEMA_signal_2953, SboxInst_n235}) ) ;
    not_masked SboxInst_U69 ( .a ({state_in_s1[97], state_in_s0[97]}), .b ({new_AGEMA_signal_2954, SboxInst_n239}) ) ;
    not_masked SboxInst_U67 ( .a ({state_in_s1[96], state_in_s0[96]}), .b ({new_AGEMA_signal_2955, SboxInst_n240}) ) ;
    not_masked SboxInst_U65 ( .a ({state_in_s1[92], state_in_s0[92]}), .b ({new_AGEMA_signal_2956, SboxInst_n227}) ) ;
    not_masked SboxInst_U63 ( .a ({state_in_s1[91], state_in_s0[91]}), .b ({new_AGEMA_signal_2957, SboxInst_n228}) ) ;
    not_masked SboxInst_U61 ( .a ({state_in_s1[94], state_in_s0[94]}), .b ({new_AGEMA_signal_2958, SboxInst_n225}) ) ;
    not_masked SboxInst_U59 ( .a ({state_in_s1[90], state_in_s0[90]}), .b ({new_AGEMA_signal_2959, SboxInst_n229}) ) ;
    not_masked SboxInst_U57 ( .a ({state_in_s1[93], state_in_s0[93]}), .b ({new_AGEMA_signal_2960, SboxInst_n226}) ) ;
    not_masked SboxInst_U55 ( .a ({state_in_s1[89], state_in_s0[89]}), .b ({new_AGEMA_signal_2961, SboxInst_n230}) ) ;
    not_masked SboxInst_U53 ( .a ({state_in_s1[88], state_in_s0[88]}), .b ({new_AGEMA_signal_2962, SboxInst_n231}) ) ;
    not_masked SboxInst_U51 ( .a ({state_in_s1[255], state_in_s0[255]}), .b ({new_AGEMA_signal_2963, SboxInst_n323}) ) ;
    not_masked SboxInst_U49 ( .a ({state_in_s1[233], state_in_s0[233]}), .b ({new_AGEMA_signal_2964, SboxInst_n376}) ) ;
    not_masked SboxInst_U47 ( .a ({state_in_s1[224], state_in_s0[224]}), .b ({new_AGEMA_signal_2965, SboxInst_n368}) ) ;
    not_masked SboxInst_U45 ( .a ({state_in_s1[254], state_in_s0[254]}), .b ({new_AGEMA_signal_2966, SboxInst_n324}) ) ;
    not_masked SboxInst_U43 ( .a ({state_in_s1[239], state_in_s0[239]}), .b ({new_AGEMA_signal_2967, SboxInst_n369}) ) ;
    not_masked SboxInst_U41 ( .a ({state_in_s1[232], state_in_s0[232]}), .b ({new_AGEMA_signal_2968, SboxInst_n377}) ) ;
    not_masked SboxInst_U39 ( .a ({state_in_s1[238], state_in_s0[238]}), .b ({new_AGEMA_signal_2969, SboxInst_n370}) ) ;
    not_masked SboxInst_U37 ( .a ({state_in_s1[247], state_in_s0[247]}), .b ({new_AGEMA_signal_2970, SboxInst_n378}) ) ;
    not_masked SboxInst_U35 ( .a ({state_in_s1[246], state_in_s0[246]}), .b ({new_AGEMA_signal_2971, SboxInst_n379}) ) ;
    not_masked SboxInst_U33 ( .a ({state_in_s1[237], state_in_s0[237]}), .b ({new_AGEMA_signal_2972, SboxInst_n371}) ) ;
    not_masked SboxInst_U31 ( .a ({state_in_s1[236], state_in_s0[236]}), .b ({new_AGEMA_signal_2973, SboxInst_n372}) ) ;
    not_masked SboxInst_U29 ( .a ({state_in_s1[245], state_in_s0[245]}), .b ({new_AGEMA_signal_2974, SboxInst_n380}) ) ;
    not_masked SboxInst_U27 ( .a ({state_in_s1[244], state_in_s0[244]}), .b ({new_AGEMA_signal_2975, SboxInst_n381}) ) ;
    not_masked SboxInst_U25 ( .a ({state_in_s1[235], state_in_s0[235]}), .b ({new_AGEMA_signal_2976, SboxInst_n374}) ) ;
    not_masked SboxInst_U23 ( .a ({state_in_s1[243], state_in_s0[243]}), .b ({new_AGEMA_signal_2977, SboxInst_n382}) ) ;
    not_masked SboxInst_U21 ( .a ({state_in_s1[234], state_in_s0[234]}), .b ({new_AGEMA_signal_2978, SboxInst_n375}) ) ;
    not_masked SboxInst_U19 ( .a ({state_in_s1[242], state_in_s0[242]}), .b ({new_AGEMA_signal_2979, SboxInst_n383}) ) ;
    not_masked SboxInst_U17 ( .a ({state_in_s1[225], state_in_s0[225]}), .b ({new_AGEMA_signal_2980, SboxInst_n367}) ) ;
    not_masked SboxInst_U15 ( .a ({state_in_s1[231], state_in_s0[231]}), .b ({new_AGEMA_signal_2981, SboxInst_n360}) ) ;
    not_masked SboxInst_U13 ( .a ({state_in_s1[230], state_in_s0[230]}), .b ({new_AGEMA_signal_2982, SboxInst_n361}) ) ;
    not_masked SboxInst_U11 ( .a ({state_in_s1[229], state_in_s0[229]}), .b ({new_AGEMA_signal_2983, SboxInst_n363}) ) ;
    not_masked SboxInst_U9 ( .a ({state_in_s1[228], state_in_s0[228]}), .b ({new_AGEMA_signal_2984, SboxInst_n364}) ) ;
    not_masked SboxInst_U7 ( .a ({state_in_s1[227], state_in_s0[227]}), .b ({new_AGEMA_signal_2985, SboxInst_n365}) ) ;
    not_masked SboxInst_U5 ( .a ({state_in_s1[241], state_in_s0[241]}), .b ({new_AGEMA_signal_2986, SboxInst_n321}) ) ;
    not_masked SboxInst_U3 ( .a ({state_in_s1[226], state_in_s0[226]}), .b ({new_AGEMA_signal_2987, SboxInst_n366}) ) ;
    not_masked SboxInst_U1 ( .a ({state_in_s1[240], state_in_s0[240]}), .b ({new_AGEMA_signal_2988, SboxInst_n322}) ) ;
    //ClockGatingController #(2) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC2 U3225 ( .a ({state_in_s1[238], state_in_s0[238]}), .b ({new_AGEMA_signal_3125, z4[22]}), .c ({new_AGEMA_signal_3295, n3405}) ) ;
    xnor_HPC2 U3226 ( .a ({state_in_s1[302], state_in_s0[302]}), .b ({new_AGEMA_signal_3295, n3405}), .c ({new_AGEMA_signal_3585, n3926}) ) ;
    xnor_HPC2 U3227 ( .a ({state_in_s1[247], state_in_s0[247]}), .b ({new_AGEMA_signal_3117, z4[15]}), .c ({new_AGEMA_signal_3296, n3487}) ) ;
    xnor_HPC2 U3228 ( .a ({state_in_s1[311], state_in_s0[311]}), .b ({new_AGEMA_signal_3296, n3487}), .c ({new_AGEMA_signal_3586, n3664}) ) ;
    xnor_HPC2 U3229 ( .a ({new_AGEMA_signal_3585, n3926}), .b ({new_AGEMA_signal_3586, n3664}), .c ({new_AGEMA_signal_3891, n3292}) ) ;
    xnor_HPC2 U3230 ( .a ({state_in_s1[192], state_in_s0[192]}), .b ({new_AGEMA_signal_3162, z4[56]}), .c ({new_AGEMA_signal_3297, n3441}) ) ;
    xnor_HPC2 U3231 ( .a ({state_in_s1[256], state_in_s0[256]}), .b ({new_AGEMA_signal_3297, n3441}), .c ({new_AGEMA_signal_3587, n3657}) ) ;
    xnor_HPC2 U3232 ( .a ({new_AGEMA_signal_3891, n3292}), .b ({new_AGEMA_signal_3587, n3657}), .c ({state_out_s1[311], state_out_s0[311]}) ) ;
    xnor_HPC2 U3233 ( .a ({state_in_s1[240], state_in_s0[240]}), .b ({new_AGEMA_signal_3173, z4[8]}), .c ({new_AGEMA_signal_3298, n3419}) ) ;
    xnor_HPC2 U3234 ( .a ({state_in_s1[304], state_in_s0[304]}), .b ({new_AGEMA_signal_3298, n3419}), .c ({new_AGEMA_signal_3588, n3663}) ) ;
    xnor_HPC2 U3235 ( .a ({state_in_s1[210], state_in_s0[210]}), .b ({new_AGEMA_signal_3147, z4[42]}), .c ({new_AGEMA_signal_3299, n3615}) ) ;
    xnor_HPC2 U3236 ( .a ({state_in_s1[274], state_in_s0[274]}), .b ({new_AGEMA_signal_3299, n3615}), .c ({new_AGEMA_signal_3589, n3661}) ) ;
    xnor_HPC2 U3237 ( .a ({new_AGEMA_signal_3588, n3663}), .b ({new_AGEMA_signal_3589, n3661}), .c ({new_AGEMA_signal_3892, n3293}) ) ;
    xnor_HPC2 U3238 ( .a ({state_in_s1[249], state_in_s0[249]}), .b ({new_AGEMA_signal_3122, z4[1]}), .c ({new_AGEMA_signal_3300, n3668}) ) ;
    xnor_HPC2 U3239 ( .a ({state_in_s1[313], state_in_s0[313]}), .b ({new_AGEMA_signal_3300, n3668}), .c ({new_AGEMA_signal_3590, n3351}) ) ;
    xnor_HPC2 U3240 ( .a ({new_AGEMA_signal_3892, n3293}), .b ({new_AGEMA_signal_3590, n3351}), .c ({state_out_s1[313], state_out_s0[313]}) ) ;
    xnor_HPC2 U3241 ( .a ({state_in_s1[241], state_in_s0[241]}), .b ({new_AGEMA_signal_3174, z4[9]}), .c ({new_AGEMA_signal_3301, n3478}) ) ;
    xnor_HPC2 U3242 ( .a ({state_in_s1[305], state_in_s0[305]}), .b ({new_AGEMA_signal_3301, n3478}), .c ({new_AGEMA_signal_3591, n3733}) ) ;
    xnor_HPC2 U3243 ( .a ({state_in_s1[211], state_in_s0[211]}), .b ({new_AGEMA_signal_3148, z4[43]}), .c ({new_AGEMA_signal_3302, n3646}) ) ;
    xnor_HPC2 U3244 ( .a ({state_in_s1[275], state_in_s0[275]}), .b ({new_AGEMA_signal_3302, n3646}), .c ({new_AGEMA_signal_3592, n3730}) ) ;
    xnor_HPC2 U3245 ( .a ({new_AGEMA_signal_3591, n3733}), .b ({new_AGEMA_signal_3592, n3730}), .c ({new_AGEMA_signal_3893, n3294}) ) ;
    xnor_HPC2 U3246 ( .a ({state_in_s1[250], state_in_s0[250]}), .b ({new_AGEMA_signal_3133, z4[2]}), .c ({new_AGEMA_signal_3303, n3706}) ) ;
    xnor_HPC2 U3247 ( .a ({state_in_s1[314], state_in_s0[314]}), .b ({new_AGEMA_signal_3303, n3706}), .c ({new_AGEMA_signal_3593, n3360}) ) ;
    xnor_HPC2 U3248 ( .a ({new_AGEMA_signal_3893, n3294}), .b ({new_AGEMA_signal_3593, n3360}), .c ({state_out_s1[314], state_out_s0[314]}) ) ;
    xnor_HPC2 U3249 ( .a ({state_in_s1[242], state_in_s0[242]}), .b ({new_AGEMA_signal_3112, z4[10]}), .c ({new_AGEMA_signal_3304, n3396}) ) ;
    xnor_HPC2 U3250 ( .a ({state_in_s1[306], state_in_s0[306]}), .b ({new_AGEMA_signal_3304, n3396}), .c ({new_AGEMA_signal_3594, n3839}) ) ;
    xnor_HPC2 U3251 ( .a ({state_in_s1[212], state_in_s0[212]}), .b ({new_AGEMA_signal_3149, z4[44]}), .c ({new_AGEMA_signal_3305, n3692}) ) ;
    xnor_HPC2 U3252 ( .a ({state_in_s1[276], state_in_s0[276]}), .b ({new_AGEMA_signal_3305, n3692}), .c ({new_AGEMA_signal_3595, n3836}) ) ;
    xnor_HPC2 U3253 ( .a ({new_AGEMA_signal_3594, n3839}), .b ({new_AGEMA_signal_3595, n3836}), .c ({new_AGEMA_signal_3894, n3295}) ) ;
    xnor_HPC2 U3254 ( .a ({state_in_s1[251], state_in_s0[251]}), .b ({new_AGEMA_signal_3144, z4[3]}), .c ({new_AGEMA_signal_3306, n3800}) ) ;
    xnor_HPC2 U3255 ( .a ({state_in_s1[315], state_in_s0[315]}), .b ({new_AGEMA_signal_3306, n3800}), .c ({new_AGEMA_signal_3596, n3391}) ) ;
    xnor_HPC2 U3256 ( .a ({new_AGEMA_signal_3894, n3295}), .b ({new_AGEMA_signal_3596, n3391}), .c ({state_out_s1[315], state_out_s0[315]}) ) ;
    xnor_HPC2 U3257 ( .a ({state_in_s1[243], state_in_s0[243]}), .b ({new_AGEMA_signal_3113, z4[11]}), .c ({new_AGEMA_signal_3307, n3438}) ) ;
    xnor_HPC2 U3258 ( .a ({state_in_s1[307], state_in_s0[307]}), .b ({new_AGEMA_signal_3307, n3438}), .c ({new_AGEMA_signal_3597, n3929}) ) ;
    xnor_HPC2 U3259 ( .a ({state_in_s1[213], state_in_s0[213]}), .b ({new_AGEMA_signal_3150, z4[45]}), .c ({new_AGEMA_signal_3308, n3783}) ) ;
    xnor_HPC2 U3260 ( .a ({state_in_s1[277], state_in_s0[277]}), .b ({new_AGEMA_signal_3308, n3783}), .c ({new_AGEMA_signal_3598, n3925}) ) ;
    xnor_HPC2 U3261 ( .a ({new_AGEMA_signal_3597, n3929}), .b ({new_AGEMA_signal_3598, n3925}), .c ({new_AGEMA_signal_3895, n3296}) ) ;
    xnor_HPC2 U3262 ( .a ({state_in_s1[252], state_in_s0[252]}), .b ({new_AGEMA_signal_3155, z4[4]}), .c ({new_AGEMA_signal_3309, n3888}) ) ;
    xnor_HPC2 U3263 ( .a ({state_in_s1[316], state_in_s0[316]}), .b ({new_AGEMA_signal_3309, n3888}), .c ({new_AGEMA_signal_3599, n3454}) ) ;
    xnor_HPC2 U3264 ( .a ({new_AGEMA_signal_3895, n3296}), .b ({new_AGEMA_signal_3599, n3454}), .c ({state_out_s1[316], state_out_s0[316]}) ) ;
    xnor_HPC2 U3265 ( .a ({state_in_s1[235], state_in_s0[235]}), .b ({new_AGEMA_signal_3121, z4[19]}), .c ({new_AGEMA_signal_3310, n3355}) ) ;
    xnor_HPC2 U3266 ( .a ({state_in_s1[299], state_in_s0[299]}), .b ({new_AGEMA_signal_3310, n3355}), .c ({new_AGEMA_signal_3600, n3660}) ) ;
    xnor_HPC2 U3267 ( .a ({state_in_s1[205], state_in_s0[205]}), .b ({new_AGEMA_signal_3159, z4[53]}), .c ({new_AGEMA_signal_3311, n3566}) ) ;
    xnor_HPC2 U3268 ( .a ({state_in_s1[269], state_in_s0[269]}), .b ({new_AGEMA_signal_3311, n3566}), .c ({new_AGEMA_signal_3601, n3625}) ) ;
    xnor_HPC2 U3269 ( .a ({new_AGEMA_signal_3600, n3660}), .b ({new_AGEMA_signal_3601, n3625}), .c ({new_AGEMA_signal_3896, n3297}) ) ;
    xnor_HPC2 U3270 ( .a ({state_in_s1[244], state_in_s0[244]}), .b ({new_AGEMA_signal_3114, z4[12]}), .c ({new_AGEMA_signal_3312, n3493}) ) ;
    xnor_HPC2 U3271 ( .a ({state_in_s1[308], state_in_s0[308]}), .b ({new_AGEMA_signal_3312, n3493}), .c ({new_AGEMA_signal_3602, n3304}) ) ;
    xnor_HPC2 U3272 ( .a ({new_AGEMA_signal_3896, n3297}), .b ({new_AGEMA_signal_3602, n3304}), .c ({state_out_s1[308], state_out_s0[308]}) ) ;
    xnor_HPC2 U3273 ( .a ({state_in_s1[214], state_in_s0[214]}), .b ({new_AGEMA_signal_3151, z4[46]}), .c ({new_AGEMA_signal_3313, n3844}) ) ;
    xnor_HPC2 U3274 ( .a ({state_in_s1[278], state_in_s0[278]}), .b ({new_AGEMA_signal_3313, n3844}), .c ({new_AGEMA_signal_3603, n3687}) ) ;
    xnor_HPC2 U3275 ( .a ({new_AGEMA_signal_3602, n3304}), .b ({new_AGEMA_signal_3603, n3687}), .c ({new_AGEMA_signal_3897, n3298}) ) ;
    xnor_HPC2 U3276 ( .a ({state_in_s1[253], state_in_s0[253]}), .b ({new_AGEMA_signal_3166, z4[5]}), .c ({new_AGEMA_signal_3314, n3738}) ) ;
    xnor_HPC2 U3277 ( .a ({state_in_s1[317], state_in_s0[317]}), .b ({new_AGEMA_signal_3314, n3738}), .c ({new_AGEMA_signal_3604, n3508}) ) ;
    xnor_HPC2 U3278 ( .a ({new_AGEMA_signal_3897, n3298}), .b ({new_AGEMA_signal_3604, n3508}), .c ({state_out_s1[317], state_out_s0[317]}) ) ;
    xnor_HPC2 U3279 ( .a ({state_in_s1[236], state_in_s0[236]}), .b ({new_AGEMA_signal_3123, z4[20]}), .c ({new_AGEMA_signal_3315, n3439}) ) ;
    xnor_HPC2 U3280 ( .a ({state_in_s1[300], state_in_s0[300]}), .b ({new_AGEMA_signal_3315, n3439}), .c ({new_AGEMA_signal_3605, n3729}) ) ;
    xnor_HPC2 U3281 ( .a ({state_in_s1[206], state_in_s0[206]}), .b ({new_AGEMA_signal_3160, z4[54]}), .c ({new_AGEMA_signal_3316, n3582}) ) ;
    xnor_HPC2 U3282 ( .a ({state_in_s1[270], state_in_s0[270]}), .b ({new_AGEMA_signal_3316, n3582}), .c ({new_AGEMA_signal_3606, n3457}) ) ;
    xnor_HPC2 U3283 ( .a ({new_AGEMA_signal_3605, n3729}), .b ({new_AGEMA_signal_3606, n3457}), .c ({new_AGEMA_signal_3898, n3299}) ) ;
    xnor_HPC2 U3284 ( .a ({state_in_s1[245], state_in_s0[245]}), .b ({new_AGEMA_signal_3115, z4[13]}), .c ({new_AGEMA_signal_3317, n3404}) ) ;
    xnor_HPC2 U3285 ( .a ({state_in_s1[309], state_in_s0[309]}), .b ({new_AGEMA_signal_3317, n3404}), .c ({new_AGEMA_signal_3607, n3306}) ) ;
    xnor_HPC2 U3286 ( .a ({new_AGEMA_signal_3898, n3299}), .b ({new_AGEMA_signal_3607, n3306}), .c ({state_out_s1[309], state_out_s0[309]}) ) ;
    xnor_HPC2 U3287 ( .a ({state_in_s1[215], state_in_s0[215]}), .b ({new_AGEMA_signal_3152, z4[47]}), .c ({new_AGEMA_signal_3318, n3354}) ) ;
    xnor_HPC2 U3288 ( .a ({state_in_s1[279], state_in_s0[279]}), .b ({new_AGEMA_signal_3318, n3354}), .c ({new_AGEMA_signal_3608, n3777}) ) ;
    xnor_HPC2 U3289 ( .a ({new_AGEMA_signal_3607, n3306}), .b ({new_AGEMA_signal_3608, n3777}), .c ({new_AGEMA_signal_3899, n3300}) ) ;
    xnor_HPC2 U3290 ( .a ({state_in_s1[254], state_in_s0[254]}), .b ({new_AGEMA_signal_3171, z4[6]}), .c ({new_AGEMA_signal_3319, n3757}) ) ;
    xnor_HPC2 U3291 ( .a ({state_in_s1[318], state_in_s0[318]}), .b ({new_AGEMA_signal_3319, n3757}), .c ({new_AGEMA_signal_3609, n3561}) ) ;
    xnor_HPC2 U3292 ( .a ({new_AGEMA_signal_3899, n3300}), .b ({new_AGEMA_signal_3609, n3561}), .c ({state_out_s1[318], state_out_s0[318]}) ) ;
    xnor_HPC2 U3293 ( .a ({state_in_s1[223], state_in_s0[223]}), .b ({new_AGEMA_signal_3143, z4[39]}), .c ({new_AGEMA_signal_3320, n3526}) ) ;
    xnor_HPC2 U3294 ( .a ({state_in_s1[287], state_in_s0[287]}), .b ({new_AGEMA_signal_3320, n3526}), .c ({new_AGEMA_signal_3610, n3686}) ) ;
    xnor_HPC2 U3295 ( .a ({new_AGEMA_signal_3591, n3733}), .b ({new_AGEMA_signal_3610, n3686}), .c ({new_AGEMA_signal_3900, n3301}) ) ;
    xnor_HPC2 U3296 ( .a ({state_in_s1[216], state_in_s0[216]}), .b ({new_AGEMA_signal_3136, z4[32]}), .c ({new_AGEMA_signal_3321, n3603}) ) ;
    xnor_HPC2 U3297 ( .a ({state_in_s1[280], state_in_s0[280]}), .b ({new_AGEMA_signal_3321, n3603}), .c ({new_AGEMA_signal_3611, n3511}) ) ;
    xnor_HPC2 U3298 ( .a ({new_AGEMA_signal_3900, n3301}), .b ({new_AGEMA_signal_3611, n3511}), .c ({state_out_s1[280], state_out_s0[280]}) ) ;
    xnor_HPC2 U3299 ( .a ({state_in_s1[208], state_in_s0[208]}), .b ({new_AGEMA_signal_3145, z4[40]}), .c ({new_AGEMA_signal_3322, n3550}) ) ;
    xnor_HPC2 U3300 ( .a ({state_in_s1[272], state_in_s0[272]}), .b ({new_AGEMA_signal_3322, n3550}), .c ({new_AGEMA_signal_3612, n3776}) ) ;
    xnor_HPC2 U3301 ( .a ({new_AGEMA_signal_3594, n3839}), .b ({new_AGEMA_signal_3612, n3776}), .c ({new_AGEMA_signal_3901, n3302}) ) ;
    xnor_HPC2 U3302 ( .a ({state_in_s1[217], state_in_s0[217]}), .b ({new_AGEMA_signal_3137, z4[33]}), .c ({new_AGEMA_signal_3323, n3613}) ) ;
    xnor_HPC2 U3303 ( .a ({state_in_s1[281], state_in_s0[281]}), .b ({new_AGEMA_signal_3323, n3613}), .c ({new_AGEMA_signal_3613, n3559}) ) ;
    xnor_HPC2 U3304 ( .a ({new_AGEMA_signal_3901, n3302}), .b ({new_AGEMA_signal_3613, n3559}), .c ({state_out_s1[281], state_out_s0[281]}) ) ;
    xnor_HPC2 U3305 ( .a ({state_in_s1[209], state_in_s0[209]}), .b ({new_AGEMA_signal_3146, z4[41]}), .c ({new_AGEMA_signal_3324, n3605}) ) ;
    xnor_HPC2 U3306 ( .a ({state_in_s1[273], state_in_s0[273]}), .b ({new_AGEMA_signal_3324, n3605}), .c ({new_AGEMA_signal_3614, n3867}) ) ;
    xnor_HPC2 U3307 ( .a ({new_AGEMA_signal_3597, n3929}), .b ({new_AGEMA_signal_3614, n3867}), .c ({new_AGEMA_signal_3902, n3303}) ) ;
    xnor_HPC2 U3308 ( .a ({state_in_s1[218], state_in_s0[218]}), .b ({new_AGEMA_signal_3138, z4[34]}), .c ({new_AGEMA_signal_3325, n3568}) ) ;
    xnor_HPC2 U3309 ( .a ({state_in_s1[282], state_in_s0[282]}), .b ({new_AGEMA_signal_3325, n3568}), .c ({new_AGEMA_signal_3615, n3422}) ) ;
    xnor_HPC2 U3310 ( .a ({new_AGEMA_signal_3902, n3303}), .b ({new_AGEMA_signal_3615, n3422}), .c ({state_out_s1[282], state_out_s0[282]}) ) ;
    xnor_HPC2 U3311 ( .a ({new_AGEMA_signal_3589, n3661}), .b ({new_AGEMA_signal_3602, n3304}), .c ({new_AGEMA_signal_3903, n3305}) ) ;
    xnor_HPC2 U3312 ( .a ({state_in_s1[219], state_in_s0[219]}), .b ({new_AGEMA_signal_3139, z4[35]}), .c ({new_AGEMA_signal_3326, n3580}) ) ;
    xnor_HPC2 U3313 ( .a ({state_in_s1[283], state_in_s0[283]}), .b ({new_AGEMA_signal_3326, n3580}), .c ({new_AGEMA_signal_3616, n3481}) ) ;
    xnor_HPC2 U3314 ( .a ({new_AGEMA_signal_3903, n3305}), .b ({new_AGEMA_signal_3616, n3481}), .c ({state_out_s1[283], state_out_s0[283]}) ) ;
    xnor_HPC2 U3315 ( .a ({new_AGEMA_signal_3592, n3730}), .b ({new_AGEMA_signal_3607, n3306}), .c ({new_AGEMA_signal_3904, n3307}) ) ;
    xnor_HPC2 U3316 ( .a ({state_in_s1[220], state_in_s0[220]}), .b ({new_AGEMA_signal_3140, z4[36]}), .c ({new_AGEMA_signal_3327, n3418}) ) ;
    xnor_HPC2 U3317 ( .a ({state_in_s1[284], state_in_s0[284]}), .b ({new_AGEMA_signal_3327, n3418}), .c ({new_AGEMA_signal_3617, n3538}) ) ;
    xnor_HPC2 U3318 ( .a ({new_AGEMA_signal_3904, n3307}), .b ({new_AGEMA_signal_3617, n3538}), .c ({state_out_s1[284], state_out_s0[284]}) ) ;
    xnor_HPC2 U3319 ( .a ({state_in_s1[221], state_in_s0[221]}), .b ({new_AGEMA_signal_3141, z4[37]}), .c ({new_AGEMA_signal_3328, n3477}) ) ;
    xnor_HPC2 U3320 ( .a ({state_in_s1[285], state_in_s0[285]}), .b ({new_AGEMA_signal_3328, n3477}), .c ({new_AGEMA_signal_3618, n3629}) ) ;
    xnor_HPC2 U3321 ( .a ({new_AGEMA_signal_3595, n3836}), .b ({new_AGEMA_signal_3618, n3629}), .c ({new_AGEMA_signal_3905, n3308}) ) ;
    xnor_HPC2 U3322 ( .a ({state_in_s1[246], state_in_s0[246]}), .b ({new_AGEMA_signal_3116, z4[14]}), .c ({new_AGEMA_signal_3329, n3598}) ) ;
    xnor_HPC2 U3323 ( .a ({state_in_s1[310], state_in_s0[310]}), .b ({new_AGEMA_signal_3329, n3598}), .c ({new_AGEMA_signal_3619, n3377}) ) ;
    xnor_HPC2 U3324 ( .a ({new_AGEMA_signal_3905, n3308}), .b ({new_AGEMA_signal_3619, n3377}), .c ({state_out_s1[285], state_out_s0[285]}) ) ;
    xnor_HPC2 U3325 ( .a ({state_in_s1[237], state_in_s0[237]}), .b ({new_AGEMA_signal_3124, z4[21]}), .c ({new_AGEMA_signal_3330, n3494}) ) ;
    xnor_HPC2 U3326 ( .a ({state_in_s1[301], state_in_s0[301]}), .b ({new_AGEMA_signal_3330, n3494}), .c ({new_AGEMA_signal_3620, n3835}) ) ;
    xnor_HPC2 U3327 ( .a ({new_AGEMA_signal_3619, n3377}), .b ({new_AGEMA_signal_3620, n3835}), .c ({new_AGEMA_signal_3906, n3309}) ) ;
    xnor_HPC2 U3328 ( .a ({state_in_s1[207], state_in_s0[207]}), .b ({new_AGEMA_signal_3161, z4[55]}), .c ({new_AGEMA_signal_3331, n3394}) ) ;
    xnor_HPC2 U3329 ( .a ({state_in_s1[271], state_in_s0[271]}), .b ({new_AGEMA_signal_3331, n3394}), .c ({new_AGEMA_signal_3621, n3510}) ) ;
    xnor_HPC2 U3330 ( .a ({new_AGEMA_signal_3906, n3309}), .b ({new_AGEMA_signal_3621, n3510}), .c ({state_out_s1[310], state_out_s0[310]}) ) ;
    xor_HPC2 U3331 ( .a ({new_AGEMA_signal_3249, z0[58]}), .b ({state_in_s1[2], state_in_s0[2]}), .c ({new_AGEMA_signal_3332, n3407}) ) ;
    xor_HPC2 U3332 ( .a ({new_AGEMA_signal_3039, z1[58]}), .b ({new_AGEMA_signal_3332, n3407}), .c ({new_AGEMA_signal_3622, n3311}) ) ;
    xnor_HPC2 U3334 ( .a ({new_AGEMA_signal_3622, n3311}), .b ({new_AGEMA_signal_2657, n3310}), .c ({new_AGEMA_signal_3907, n3542}) ) ;
    xor_HPC2 U3335 ( .a ({new_AGEMA_signal_3014, z1[33]}), .b ({state_in_s1[281], state_in_s0[281]}), .c ({new_AGEMA_signal_3333, n3313}) ) ;
    xor_HPC2 U3336 ( .a ({new_AGEMA_signal_3267, z0[33]}), .b ({state_in_s1[25], state_in_s0[25]}), .c ({new_AGEMA_signal_3334, n3614}) ) ;
    xnor_HPC2 U3337 ( .a ({state_in_s1[89], state_in_s0[89]}), .b ({new_AGEMA_signal_3334, n3614}), .c ({new_AGEMA_signal_3623, n3312}) ) ;
    xnor_HPC2 U3338 ( .a ({new_AGEMA_signal_3333, n3313}), .b ({new_AGEMA_signal_3623, n3312}), .c ({new_AGEMA_signal_3908, n3447}) ) ;
    xnor_HPC2 U3339 ( .a ({new_AGEMA_signal_3907, n3542}), .b ({new_AGEMA_signal_3908, n3447}), .c ({new_AGEMA_signal_4220, n3316}) ) ;
    xor_HPC2 U3340 ( .a ({new_AGEMA_signal_3036, z1[55]}), .b ({state_in_s1[271], state_in_s0[271]}), .c ({new_AGEMA_signal_3335, n3315}) ) ;
    xor_HPC2 U3341 ( .a ({new_AGEMA_signal_3253, z0[55]}), .b ({state_in_s1[15], state_in_s0[15]}), .c ({new_AGEMA_signal_3336, n3395}) ) ;
    xnor_HPC2 U3342 ( .a ({state_in_s1[79], state_in_s0[79]}), .b ({new_AGEMA_signal_3336, n3395}), .c ({new_AGEMA_signal_3624, n3314}) ) ;
    xnor_HPC2 U3343 ( .a ({new_AGEMA_signal_3335, n3315}), .b ({new_AGEMA_signal_3624, n3314}), .c ({new_AGEMA_signal_3909, n3433}) ) ;
    xnor_HPC2 U3344 ( .a ({new_AGEMA_signal_4220, n3316}), .b ({new_AGEMA_signal_3909, n3433}), .c ({state_out_s1[66], state_out_s0[66]}) ) ;
    xor_HPC2 U3345 ( .a ({new_AGEMA_signal_3247, z0[59]}), .b ({state_in_s1[3], state_in_s0[3]}), .c ({new_AGEMA_signal_3337, n3597}) ) ;
    xor_HPC2 U3346 ( .a ({new_AGEMA_signal_3040, z1[59]}), .b ({new_AGEMA_signal_3337, n3597}), .c ({new_AGEMA_signal_3625, n3318}) ) ;
    xnor_HPC2 U3348 ( .a ({new_AGEMA_signal_3625, n3318}), .b ({new_AGEMA_signal_2659, n3317}), .c ({new_AGEMA_signal_3910, n3572}) ) ;
    xor_HPC2 U3349 ( .a ({new_AGEMA_signal_3015, z1[34]}), .b ({state_in_s1[282], state_in_s0[282]}), .c ({new_AGEMA_signal_3338, n3320}) ) ;
    xor_HPC2 U3350 ( .a ({new_AGEMA_signal_3265, z0[34]}), .b ({state_in_s1[26], state_in_s0[26]}), .c ({new_AGEMA_signal_3339, n3569}) ) ;
    xnor_HPC2 U3351 ( .a ({state_in_s1[90], state_in_s0[90]}), .b ({new_AGEMA_signal_3339, n3569}), .c ({new_AGEMA_signal_3626, n3319}) ) ;
    xnor_HPC2 U3352 ( .a ({new_AGEMA_signal_3338, n3320}), .b ({new_AGEMA_signal_3626, n3319}), .c ({new_AGEMA_signal_3911, n3502}) ) ;
    xnor_HPC2 U3353 ( .a ({new_AGEMA_signal_3910, n3572}), .b ({new_AGEMA_signal_3911, n3502}), .c ({new_AGEMA_signal_4221, n3323}) ) ;
    xor_HPC2 U3354 ( .a ({new_AGEMA_signal_3037, z1[56]}), .b ({state_in_s1[256], state_in_s0[256]}), .c ({new_AGEMA_signal_3340, n3322}) ) ;
    xor_HPC2 U3355 ( .a ({new_AGEMA_signal_3252, z0[56]}), .b ({state_in_s1[0], state_in_s0[0]}), .c ({new_AGEMA_signal_3341, n3442}) ) ;
    xnor_HPC2 U3356 ( .a ({state_in_s1[64], state_in_s0[64]}), .b ({new_AGEMA_signal_3341, n3442}), .c ({new_AGEMA_signal_3627, n3321}) ) ;
    xnor_HPC2 U3357 ( .a ({new_AGEMA_signal_3340, n3322}), .b ({new_AGEMA_signal_3627, n3321}), .c ({new_AGEMA_signal_3912, n3464}) ) ;
    xnor_HPC2 U3358 ( .a ({new_AGEMA_signal_4221, n3323}), .b ({new_AGEMA_signal_3912, n3464}), .c ({state_out_s1[67], state_out_s0[67]}) ) ;
    xnor_HPC2 U3359 ( .a ({new_AGEMA_signal_3586, n3664}), .b ({new_AGEMA_signal_3598, n3925}), .c ({new_AGEMA_signal_3913, n3324}) ) ;
    xnor_HPC2 U3360 ( .a ({state_in_s1[222], state_in_s0[222]}), .b ({new_AGEMA_signal_3142, z4[38]}), .c ({new_AGEMA_signal_3342, n3353}) ) ;
    xnor_HPC2 U3361 ( .a ({state_in_s1[286], state_in_s0[286]}), .b ({new_AGEMA_signal_3342, n3353}), .c ({new_AGEMA_signal_3628, n3453}) ) ;
    xnor_HPC2 U3362 ( .a ({new_AGEMA_signal_3913, n3324}), .b ({new_AGEMA_signal_3628, n3453}), .c ({state_out_s1[286], state_out_s0[286]}) ) ;
    xnor_HPC2 U3363 ( .a ({new_AGEMA_signal_3588, n3663}), .b ({new_AGEMA_signal_3628, n3453}), .c ({new_AGEMA_signal_3914, n3325}) ) ;
    xnor_HPC2 U3364 ( .a ({state_in_s1[231], state_in_s0[231]}), .b ({new_AGEMA_signal_3135, z4[31]}), .c ({new_AGEMA_signal_3343, n3551}) ) ;
    xnor_HPC2 U3365 ( .a ({state_in_s1[295], state_in_s0[295]}), .b ({new_AGEMA_signal_3343, n3551}), .c ({new_AGEMA_signal_3629, n3456}) ) ;
    xnor_HPC2 U3366 ( .a ({new_AGEMA_signal_3914, n3325}), .b ({new_AGEMA_signal_3629, n3456}), .c ({state_out_s1[295], state_out_s0[295]}) ) ;
    xnor_HPC2 U3367 ( .a ({state_in_s1[193], state_in_s0[193]}), .b ({new_AGEMA_signal_3163, z4[57]}), .c ({new_AGEMA_signal_3344, n3496}) ) ;
    xnor_HPC2 U3368 ( .a ({state_in_s1[257], state_in_s0[257]}), .b ({new_AGEMA_signal_3344, n3496}), .c ({new_AGEMA_signal_3630, n3726}) ) ;
    xnor_HPC2 U3369 ( .a ({new_AGEMA_signal_3615, n3422}), .b ({new_AGEMA_signal_3630, n3726}), .c ({new_AGEMA_signal_3915, n3326}) ) ;
    xnor_HPC2 U3370 ( .a ({state_in_s1[248], state_in_s0[248]}), .b ({new_AGEMA_signal_3111, z4[0]}), .c ({new_AGEMA_signal_3345, n3634}) ) ;
    xnor_HPC2 U3371 ( .a ({state_in_s1[312], state_in_s0[312]}), .b ({new_AGEMA_signal_3345, n3634}), .c ({new_AGEMA_signal_3631, n3631}) ) ;
    xnor_HPC2 U3372 ( .a ({new_AGEMA_signal_3915, n3326}), .b ({new_AGEMA_signal_3631, n3631}), .c ({state_out_s1[257], state_out_s0[257]}) ) ;
    xor_HPC2 U3373 ( .a ({new_AGEMA_signal_3041, z1[60]}), .b ({state_in_s1[260], state_in_s0[260]}), .c ({new_AGEMA_signal_3346, n3328}) ) ;
    xor_HPC2 U3374 ( .a ({new_AGEMA_signal_3244, z0[60]}), .b ({state_in_s1[4], state_in_s0[4]}), .c ({new_AGEMA_signal_3347, n3486}) ) ;
    xnor_HPC2 U3375 ( .a ({state_in_s1[68], state_in_s0[68]}), .b ({new_AGEMA_signal_3347, n3486}), .c ({new_AGEMA_signal_3632, n3327}) ) ;
    xnor_HPC2 U3376 ( .a ({new_AGEMA_signal_3346, n3328}), .b ({new_AGEMA_signal_3632, n3327}), .c ({new_AGEMA_signal_3916, n3586}) ) ;
    xor_HPC2 U3377 ( .a ({new_AGEMA_signal_3251, z0[57]}), .b ({state_in_s1[1], state_in_s0[1]}), .c ({new_AGEMA_signal_3348, n3497}) ) ;
    xor_HPC2 U3378 ( .a ({new_AGEMA_signal_3038, z1[57]}), .b ({new_AGEMA_signal_3348, n3497}), .c ({new_AGEMA_signal_3633, n3330}) ) ;
    xnor_HPC2 U3380 ( .a ({new_AGEMA_signal_3633, n3330}), .b ({new_AGEMA_signal_2661, n3329}), .c ({new_AGEMA_signal_3917, n3515}) ) ;
    xnor_HPC2 U3381 ( .a ({new_AGEMA_signal_3916, n3586}), .b ({new_AGEMA_signal_3917, n3515}), .c ({new_AGEMA_signal_4225, n3333}) ) ;
    xor_HPC2 U3382 ( .a ({new_AGEMA_signal_3016, z1[35]}), .b ({state_in_s1[283], state_in_s0[283]}), .c ({new_AGEMA_signal_3349, n3332}) ) ;
    xor_HPC2 U3383 ( .a ({new_AGEMA_signal_3263, z0[35]}), .b ({state_in_s1[27], state_in_s0[27]}), .c ({new_AGEMA_signal_3350, n3581}) ) ;
    xnor_HPC2 U3384 ( .a ({state_in_s1[91], state_in_s0[91]}), .b ({new_AGEMA_signal_3350, n3581}), .c ({new_AGEMA_signal_3634, n3331}) ) ;
    xnor_HPC2 U3385 ( .a ({new_AGEMA_signal_3349, n3332}), .b ({new_AGEMA_signal_3634, n3331}), .c ({new_AGEMA_signal_3918, n3412}) ) ;
    xnor_HPC2 U3386 ( .a ({new_AGEMA_signal_4225, n3333}), .b ({new_AGEMA_signal_3918, n3412}), .c ({state_out_s1[68], state_out_s0[68]}) ) ;
    xor_HPC2 U3387 ( .a ({new_AGEMA_signal_3002, z1[21]}), .b ({state_in_s1[301], state_in_s0[301]}), .c ({new_AGEMA_signal_3351, n3335}) ) ;
    xor_HPC2 U3388 ( .a ({new_AGEMA_signal_3245, z0[21]}), .b ({state_in_s1[45], state_in_s0[45]}), .c ({new_AGEMA_signal_3352, n3495}) ) ;
    xnor_HPC2 U3389 ( .a ({state_in_s1[109], state_in_s0[109]}), .b ({new_AGEMA_signal_3352, n3495}), .c ({new_AGEMA_signal_3635, n3334}) ) ;
    xnor_HPC2 U3390 ( .a ({new_AGEMA_signal_3351, n3335}), .b ({new_AGEMA_signal_3635, n3334}), .c ({new_AGEMA_signal_3919, n3853}) ) ;
    xnor_HPC2 U3391 ( .a ({new_AGEMA_signal_3916, n3586}), .b ({new_AGEMA_signal_3919, n3853}), .c ({new_AGEMA_signal_4226, n3338}) ) ;
    xor_HPC2 U3392 ( .a ({new_AGEMA_signal_3246, z0[18]}), .b ({state_in_s1[42], state_in_s0[42]}), .c ({new_AGEMA_signal_3353, n3857}) ) ;
    xor_HPC2 U3393 ( .a ({new_AGEMA_signal_2999, z1[18]}), .b ({new_AGEMA_signal_3353, n3857}), .c ({new_AGEMA_signal_3636, n3337}) ) ;
    xnor_HPC2 U3395 ( .a ({new_AGEMA_signal_3636, n3337}), .b ({new_AGEMA_signal_2663, n3336}), .c ({new_AGEMA_signal_3920, n3648}) ) ;
    xnor_HPC2 U3396 ( .a ({new_AGEMA_signal_4226, n3338}), .b ({new_AGEMA_signal_3920, n3648}), .c ({state_out_s1[109], state_out_s0[109]}) ) ;
    xor_HPC2 U3397 ( .a ({new_AGEMA_signal_3000, z1[19]}), .b ({state_in_s1[299], state_in_s0[299]}), .c ({new_AGEMA_signal_3354, n3340}) ) ;
    xor_HPC2 U3398 ( .a ({new_AGEMA_signal_3242, z0[19]}), .b ({state_in_s1[43], state_in_s0[43]}), .c ({new_AGEMA_signal_3355, n3356}) ) ;
    xnor_HPC2 U3399 ( .a ({state_in_s1[107], state_in_s0[107]}), .b ({new_AGEMA_signal_3355, n3356}), .c ({new_AGEMA_signal_3637, n3339}) ) ;
    xnor_HPC2 U3400 ( .a ({new_AGEMA_signal_3354, n3340}), .b ({new_AGEMA_signal_3637, n3339}), .c ({new_AGEMA_signal_3921, n3697}) ) ;
    xnor_HPC2 U3401 ( .a ({new_AGEMA_signal_3907, n3542}), .b ({new_AGEMA_signal_3921, n3697}), .c ({new_AGEMA_signal_4227, n3343}) ) ;
    xor_HPC2 U3402 ( .a ({new_AGEMA_signal_2997, z1[16]}), .b ({state_in_s1[296], state_in_s0[296]}), .c ({new_AGEMA_signal_3356, n3342}) ) ;
    xor_HPC2 U3403 ( .a ({new_AGEMA_signal_3250, z0[16]}), .b ({state_in_s1[40], state_in_s0[40]}), .c ({new_AGEMA_signal_3357, n3682}) ) ;
    xnor_HPC2 U3404 ( .a ({state_in_s1[104], state_in_s0[104]}), .b ({new_AGEMA_signal_3357, n3682}), .c ({new_AGEMA_signal_3638, n3341}) ) ;
    xnor_HPC2 U3405 ( .a ({new_AGEMA_signal_3356, n3342}), .b ({new_AGEMA_signal_3638, n3341}), .c ({new_AGEMA_signal_3922, n3608}) ) ;
    xnor_HPC2 U3406 ( .a ({new_AGEMA_signal_4227, n3343}), .b ({new_AGEMA_signal_3922, n3608}), .c ({state_out_s1[107], state_out_s0[107]}) ) ;
    xnor_HPC2 U3407 ( .a ({new_AGEMA_signal_3606, n3457}), .b ({new_AGEMA_signal_3608, n3777}), .c ({new_AGEMA_signal_3923, n3344}) ) ;
    xnor_HPC2 U3408 ( .a ({state_in_s1[224], state_in_s0[224]}), .b ({new_AGEMA_signal_3127, z4[24]}), .c ({new_AGEMA_signal_3358, n3484}) ) ;
    xnor_HPC2 U3409 ( .a ({state_in_s1[288], state_in_s0[288]}), .b ({new_AGEMA_signal_3358, n3484}), .c ({new_AGEMA_signal_3639, n3780}) ) ;
    xnor_HPC2 U3410 ( .a ({new_AGEMA_signal_3923, n3344}), .b ({new_AGEMA_signal_3639, n3780}), .c ({state_out_s1[279], state_out_s0[279]}) ) ;
    xnor_HPC2 U3411 ( .a ({new_AGEMA_signal_3590, n3351}), .b ({new_AGEMA_signal_3629, n3456}), .c ({new_AGEMA_signal_3924, n3345}) ) ;
    xnor_HPC2 U3412 ( .a ({new_AGEMA_signal_3924, n3345}), .b ({new_AGEMA_signal_3639, n3780}), .c ({state_out_s1[288], state_out_s0[288]}) ) ;
    xor_HPC2 U3413 ( .a ({new_AGEMA_signal_3001, z1[20]}), .b ({state_in_s1[300], state_in_s0[300]}), .c ({new_AGEMA_signal_3359, n3347}) ) ;
    xor_HPC2 U3414 ( .a ({new_AGEMA_signal_3240, z0[20]}), .b ({state_in_s1[44], state_in_s0[44]}), .c ({new_AGEMA_signal_3360, n3440}) ) ;
    xnor_HPC2 U3415 ( .a ({state_in_s1[108], state_in_s0[108]}), .b ({new_AGEMA_signal_3360, n3440}), .c ({new_AGEMA_signal_3640, n3346}) ) ;
    xnor_HPC2 U3416 ( .a ({new_AGEMA_signal_3359, n3347}), .b ({new_AGEMA_signal_3640, n3346}), .c ({new_AGEMA_signal_3925, n3796}) ) ;
    xnor_HPC2 U3417 ( .a ({new_AGEMA_signal_3910, n3572}), .b ({new_AGEMA_signal_3925, n3796}), .c ({new_AGEMA_signal_4230, n3350}) ) ;
    xor_HPC2 U3418 ( .a ({new_AGEMA_signal_3248, z0[17]}), .b ({state_in_s1[41], state_in_s0[41]}), .c ({new_AGEMA_signal_3361, n3771}) ) ;
    xor_HPC2 U3419 ( .a ({new_AGEMA_signal_2998, z1[17]}), .b ({new_AGEMA_signal_3361, n3771}), .c ({new_AGEMA_signal_3641, n3349}) ) ;
    xnor_HPC2 U3421 ( .a ({new_AGEMA_signal_3641, n3349}), .b ({new_AGEMA_signal_2665, n3348}), .c ({new_AGEMA_signal_3926, n3617}) ) ;
    xnor_HPC2 U3422 ( .a ({new_AGEMA_signal_4230, n3350}), .b ({new_AGEMA_signal_3926, n3617}), .c ({state_out_s1[108], state_out_s0[108]}) ) ;
    xnor_HPC2 U3423 ( .a ({new_AGEMA_signal_3590, n3351}), .b ({new_AGEMA_signal_3616, n3481}), .c ({new_AGEMA_signal_3927, n3352}) ) ;
    xnor_HPC2 U3424 ( .a ({state_in_s1[194], state_in_s0[194]}), .b ({new_AGEMA_signal_3164, z4[58]}), .c ({new_AGEMA_signal_3362, n3406}) ) ;
    xnor_HPC2 U3425 ( .a ({state_in_s1[258], state_in_s0[258]}), .b ({new_AGEMA_signal_3362, n3406}), .c ({new_AGEMA_signal_3642, n3832}) ) ;
    xnor_HPC2 U3426 ( .a ({new_AGEMA_signal_3927, n3352}), .b ({new_AGEMA_signal_3642, n3832}), .c ({state_out_s1[258], state_out_s0[258]}) ) ;
    xor_HPC2 U3427 ( .a ({new_AGEMA_signal_3264, z0[38]}), .b ({state_in_s1[30], state_in_s0[30]}), .c ({new_AGEMA_signal_3363, n3409}) ) ;
    xnor_HPC2 U3428 ( .a ({new_AGEMA_signal_3363, n3409}), .b ({new_AGEMA_signal_3342, n3353}), .c ({new_AGEMA_signal_3643, n3709}) ) ;
    xor_HPC2 U3429 ( .a ({new_AGEMA_signal_3239, z0[47]}), .b ({state_in_s1[23], state_in_s0[23]}), .c ({new_AGEMA_signal_3364, n3369}) ) ;
    xnor_HPC2 U3430 ( .a ({new_AGEMA_signal_3364, n3369}), .b ({new_AGEMA_signal_3318, n3354}), .c ({new_AGEMA_signal_3644, n3705}) ) ;
    xnor_HPC2 U3431 ( .a ({new_AGEMA_signal_3643, n3709}), .b ({new_AGEMA_signal_3644, n3705}), .c ({new_AGEMA_signal_3928, n3357}) ) ;
    xnor_HPC2 U3432 ( .a ({new_AGEMA_signal_3355, n3356}), .b ({new_AGEMA_signal_3310, n3355}), .c ({new_AGEMA_signal_3645, n3637}) ) ;
    xnor_HPC2 U3433 ( .a ({new_AGEMA_signal_3928, n3357}), .b ({new_AGEMA_signal_3645, n3637}), .c ({state_out_s1[43], state_out_s0[43]}) ) ;
    xnor_HPC2 U3434 ( .a ({state_in_s1[225], state_in_s0[225]}), .b ({new_AGEMA_signal_3128, z4[25]}), .c ({new_AGEMA_signal_3365, n3683}) ) ;
    xnor_HPC2 U3435 ( .a ({state_in_s1[289], state_in_s0[289]}), .b ({new_AGEMA_signal_3365, n3683}), .c ({new_AGEMA_signal_3646, n3870}) ) ;
    xnor_HPC2 U3436 ( .a ({new_AGEMA_signal_3621, n3510}), .b ({new_AGEMA_signal_3646, n3870}), .c ({new_AGEMA_signal_3929, n3358}) ) ;
    xnor_HPC2 U3437 ( .a ({state_in_s1[200], state_in_s0[200]}), .b ({new_AGEMA_signal_3153, z4[48]}), .c ({new_AGEMA_signal_3366, n3527}) ) ;
    xnor_HPC2 U3438 ( .a ({state_in_s1[264], state_in_s0[264]}), .b ({new_AGEMA_signal_3366, n3527}), .c ({new_AGEMA_signal_3647, n3866}) ) ;
    xnor_HPC2 U3439 ( .a ({new_AGEMA_signal_3929, n3358}), .b ({new_AGEMA_signal_3647, n3866}), .c ({state_out_s1[264], state_out_s0[264]}) ) ;
    xnor_HPC2 U3440 ( .a ({new_AGEMA_signal_3593, n3360}), .b ({new_AGEMA_signal_3611, n3511}), .c ({new_AGEMA_signal_3930, n3359}) ) ;
    xnor_HPC2 U3441 ( .a ({new_AGEMA_signal_3930, n3359}), .b ({new_AGEMA_signal_3646, n3870}), .c ({state_out_s1[289], state_out_s0[289]}) ) ;
    xnor_HPC2 U3442 ( .a ({new_AGEMA_signal_3593, n3360}), .b ({new_AGEMA_signal_3617, n3538}), .c ({new_AGEMA_signal_3931, n3361}) ) ;
    xnor_HPC2 U3443 ( .a ({state_in_s1[195], state_in_s0[195]}), .b ({new_AGEMA_signal_3165, z4[59]}), .c ({new_AGEMA_signal_3367, n3596}) ) ;
    xnor_HPC2 U3444 ( .a ({state_in_s1[259], state_in_s0[259]}), .b ({new_AGEMA_signal_3367, n3596}), .c ({new_AGEMA_signal_3648, n3922}) ) ;
    xnor_HPC2 U3445 ( .a ({new_AGEMA_signal_3931, n3361}), .b ({new_AGEMA_signal_3648, n3922}), .c ({state_out_s1[259], state_out_s0[259]}) ) ;
    xor_HPC2 U3446 ( .a ({new_AGEMA_signal_3045, z1[8]}), .b ({state_in_s1[304], state_in_s0[304]}), .c ({new_AGEMA_signal_3368, n3363}) ) ;
    xor_HPC2 U3447 ( .a ({new_AGEMA_signal_3235, z0[8]}), .b ({state_in_s1[48], state_in_s0[48]}), .c ({new_AGEMA_signal_3369, n3420}) ) ;
    xnor_HPC2 U3448 ( .a ({state_in_s1[112], state_in_s0[112]}), .b ({new_AGEMA_signal_3369, n3420}), .c ({new_AGEMA_signal_3649, n3362}) ) ;
    xnor_HPC2 U3449 ( .a ({new_AGEMA_signal_3368, n3363}), .b ({new_AGEMA_signal_3649, n3362}), .c ({new_AGEMA_signal_3932, n3751}) ) ;
    xnor_HPC2 U3450 ( .a ({new_AGEMA_signal_3908, n3447}), .b ({new_AGEMA_signal_3932, n3751}), .c ({new_AGEMA_signal_4236, n3366}) ) ;
    xor_HPC2 U3451 ( .a ({new_AGEMA_signal_3011, z1[30]}), .b ({state_in_s1[294], state_in_s0[294]}), .c ({new_AGEMA_signal_3370, n3365}) ) ;
    xor_HPC2 U3452 ( .a ({new_AGEMA_signal_3256, z0[30]}), .b ({state_in_s1[38], state_in_s0[38]}), .c ({new_AGEMA_signal_3371, n3622}) ) ;
    xnor_HPC2 U3453 ( .a ({state_in_s1[102], state_in_s0[102]}), .b ({new_AGEMA_signal_3371, n3622}), .c ({new_AGEMA_signal_3650, n3364}) ) ;
    xnor_HPC2 U3454 ( .a ({new_AGEMA_signal_3370, n3365}), .b ({new_AGEMA_signal_3650, n3364}), .c ({new_AGEMA_signal_3933, n3745}) ) ;
    xnor_HPC2 U3455 ( .a ({new_AGEMA_signal_4236, n3366}), .b ({new_AGEMA_signal_3933, n3745}), .c ({state_out_s1[89], state_out_s0[89]}) ) ;
    xor_HPC2 U3456 ( .a ({new_AGEMA_signal_3260, z0[25]}), .b ({state_in_s1[33], state_in_s0[33]}), .c ({new_AGEMA_signal_3372, n3684}) ) ;
    xor_HPC2 U3457 ( .a ({new_AGEMA_signal_3006, z1[25]}), .b ({new_AGEMA_signal_3372, n3684}), .c ({new_AGEMA_signal_3651, n3368}) ) ;
    xnor_HPC2 U3459 ( .a ({new_AGEMA_signal_3651, n3368}), .b ({new_AGEMA_signal_2667, n3367}), .c ({new_AGEMA_signal_3934, n3810}) ) ;
    xor_HPC2 U3460 ( .a ({new_AGEMA_signal_3028, z1[47]}), .b ({new_AGEMA_signal_3364, n3369}), .c ({new_AGEMA_signal_3652, n3371}) ) ;
    xnor_HPC2 U3462 ( .a ({new_AGEMA_signal_3652, n3371}), .b ({new_AGEMA_signal_2669, n3370}), .c ({new_AGEMA_signal_3935, n3750}) ) ;
    xnor_HPC2 U3463 ( .a ({new_AGEMA_signal_3934, n3810}), .b ({new_AGEMA_signal_3935, n3750}), .c ({new_AGEMA_signal_4237, n3374}) ) ;
    xor_HPC2 U3464 ( .a ({new_AGEMA_signal_3031, z1[50]}), .b ({state_in_s1[266], state_in_s0[266]}), .c ({new_AGEMA_signal_3373, n3373}) ) ;
    xor_HPC2 U3465 ( .a ({new_AGEMA_signal_3236, z0[50]}), .b ({state_in_s1[10], state_in_s0[10]}), .c ({new_AGEMA_signal_3374, n3722}) ) ;
    xnor_HPC2 U3466 ( .a ({state_in_s1[74], state_in_s0[74]}), .b ({new_AGEMA_signal_3374, n3722}), .c ({new_AGEMA_signal_3653, n3372}) ) ;
    xnor_HPC2 U3467 ( .a ({new_AGEMA_signal_3373, n3373}), .b ({new_AGEMA_signal_3653, n3372}), .c ({new_AGEMA_signal_3936, n3468}) ) ;
    xnor_HPC2 U3468 ( .a ({new_AGEMA_signal_4237, n3374}), .b ({new_AGEMA_signal_3936, n3468}), .c ({state_out_s1[74], state_out_s0[74]}) ) ;
    xnor_HPC2 U3469 ( .a ({new_AGEMA_signal_3596, n3391}), .b ({new_AGEMA_signal_3613, n3559}), .c ({new_AGEMA_signal_3937, n3375}) ) ;
    xnor_HPC2 U3470 ( .a ({state_in_s1[226], state_in_s0[226]}), .b ({new_AGEMA_signal_3129, z4[26]}), .c ({new_AGEMA_signal_3375, n3769}) ) ;
    xnor_HPC2 U3471 ( .a ({state_in_s1[290], state_in_s0[290]}), .b ({new_AGEMA_signal_3375, n3769}), .c ({new_AGEMA_signal_3654, n3656}) ) ;
    xnor_HPC2 U3472 ( .a ({new_AGEMA_signal_3937, n3375}), .b ({new_AGEMA_signal_3654, n3656}), .c ({state_out_s1[290], state_out_s0[290]}) ) ;
    xnor_HPC2 U3473 ( .a ({new_AGEMA_signal_3614, n3867}), .b ({new_AGEMA_signal_3631, n3631}), .c ({new_AGEMA_signal_3938, n3376}) ) ;
    xnor_HPC2 U3474 ( .a ({state_in_s1[255], state_in_s0[255]}), .b ({new_AGEMA_signal_3172, z4[7]}), .c ({new_AGEMA_signal_3376, n3873}) ) ;
    xnor_HPC2 U3475 ( .a ({state_in_s1[319], state_in_s0[319]}), .b ({new_AGEMA_signal_3376, n3873}), .c ({new_AGEMA_signal_3655, n3628}) ) ;
    xnor_HPC2 U3476 ( .a ({new_AGEMA_signal_3938, n3376}), .b ({new_AGEMA_signal_3655, n3628}), .c ({state_out_s1[312], state_out_s0[312]}) ) ;
    xnor_HPC2 U3477 ( .a ({new_AGEMA_signal_3619, n3377}), .b ({new_AGEMA_signal_3647, n3866}), .c ({new_AGEMA_signal_3939, n3378}) ) ;
    xnor_HPC2 U3478 ( .a ({new_AGEMA_signal_3939, n3378}), .b ({new_AGEMA_signal_3655, n3628}), .c ({state_out_s1[319], state_out_s0[319]}) ) ;
    xor_HPC2 U3479 ( .a ({new_AGEMA_signal_3046, z1[9]}), .b ({state_in_s1[305], state_in_s0[305]}), .c ({new_AGEMA_signal_3377, n3380}) ) ;
    xor_HPC2 U3480 ( .a ({new_AGEMA_signal_3233, z0[9]}), .b ({state_in_s1[49], state_in_s0[49]}), .c ({new_AGEMA_signal_3378, n3479}) ) ;
    xnor_HPC2 U3481 ( .a ({state_in_s1[113], state_in_s0[113]}), .b ({new_AGEMA_signal_3378, n3479}), .c ({new_AGEMA_signal_3656, n3379}) ) ;
    xnor_HPC2 U3482 ( .a ({new_AGEMA_signal_3377, n3380}), .b ({new_AGEMA_signal_3656, n3379}), .c ({new_AGEMA_signal_3940, n3767}) ) ;
    xnor_HPC2 U3483 ( .a ({new_AGEMA_signal_3911, n3502}), .b ({new_AGEMA_signal_3940, n3767}), .c ({new_AGEMA_signal_4241, n3383}) ) ;
    xor_HPC2 U3484 ( .a ({new_AGEMA_signal_3012, z1[31]}), .b ({state_in_s1[295], state_in_s0[295]}), .c ({new_AGEMA_signal_3379, n3382}) ) ;
    xor_HPC2 U3485 ( .a ({new_AGEMA_signal_3254, z0[31]}), .b ({state_in_s1[39], state_in_s0[39]}), .c ({new_AGEMA_signal_3380, n3552}) ) ;
    xnor_HPC2 U3486 ( .a ({state_in_s1[103], state_in_s0[103]}), .b ({new_AGEMA_signal_3380, n3552}), .c ({new_AGEMA_signal_3657, n3381}) ) ;
    xnor_HPC2 U3487 ( .a ({new_AGEMA_signal_3379, n3382}), .b ({new_AGEMA_signal_3657, n3381}), .c ({new_AGEMA_signal_3941, n3762}) ) ;
    xnor_HPC2 U3488 ( .a ({new_AGEMA_signal_4241, n3383}), .b ({new_AGEMA_signal_3941, n3762}), .c ({state_out_s1[90], state_out_s0[90]}) ) ;
    xor_HPC2 U3489 ( .a ({new_AGEMA_signal_3007, z1[26]}), .b ({state_in_s1[290], state_in_s0[290]}), .c ({new_AGEMA_signal_3381, n3385}) ) ;
    xor_HPC2 U3490 ( .a ({new_AGEMA_signal_3258, z0[26]}), .b ({state_in_s1[34], state_in_s0[34]}), .c ({new_AGEMA_signal_3382, n3770}) ) ;
    xnor_HPC2 U3491 ( .a ({state_in_s1[98], state_in_s0[98]}), .b ({new_AGEMA_signal_3382, n3770}), .c ({new_AGEMA_signal_3658, n3384}) ) ;
    xnor_HPC2 U3492 ( .a ({new_AGEMA_signal_3381, n3385}), .b ({new_AGEMA_signal_3658, n3384}), .c ({new_AGEMA_signal_3942, n3898}) ) ;
    xor_HPC2 U3493 ( .a ({new_AGEMA_signal_3238, z0[48]}), .b ({state_in_s1[8], state_in_s0[8]}), .c ({new_AGEMA_signal_3383, n3528}) ) ;
    xor_HPC2 U3494 ( .a ({new_AGEMA_signal_3029, z1[48]}), .b ({new_AGEMA_signal_3383, n3528}), .c ({new_AGEMA_signal_3659, n3387}) ) ;
    xnor_HPC2 U3496 ( .a ({new_AGEMA_signal_3659, n3387}), .b ({new_AGEMA_signal_2671, n3386}), .c ({new_AGEMA_signal_3943, n3791}) ) ;
    xnor_HPC2 U3497 ( .a ({new_AGEMA_signal_3942, n3898}), .b ({new_AGEMA_signal_3943, n3791}), .c ({new_AGEMA_signal_4242, n3390}) ) ;
    xor_HPC2 U3498 ( .a ({new_AGEMA_signal_3234, z0[51]}), .b ({state_in_s1[11], state_in_s0[11]}), .c ({new_AGEMA_signal_3384, n3824}) ) ;
    xor_HPC2 U3499 ( .a ({new_AGEMA_signal_3032, z1[51]}), .b ({new_AGEMA_signal_3384, n3824}), .c ({new_AGEMA_signal_3660, n3389}) ) ;
    xnor_HPC2 U3501 ( .a ({new_AGEMA_signal_3660, n3389}), .b ({new_AGEMA_signal_2673, n3388}), .c ({new_AGEMA_signal_3944, n3519}) ) ;
    xnor_HPC2 U3502 ( .a ({new_AGEMA_signal_4242, n3390}), .b ({new_AGEMA_signal_3944, n3519}), .c ({state_out_s1[75], state_out_s0[75]}) ) ;
    xnor_HPC2 U3503 ( .a ({new_AGEMA_signal_3596, n3391}), .b ({new_AGEMA_signal_3618, n3629}), .c ({new_AGEMA_signal_3945, n3392}) ) ;
    xnor_HPC2 U3504 ( .a ({state_in_s1[196], state_in_s0[196]}), .b ({new_AGEMA_signal_3167, z4[60]}), .c ({new_AGEMA_signal_3385, n3485}) ) ;
    xnor_HPC2 U3505 ( .a ({state_in_s1[260], state_in_s0[260]}), .b ({new_AGEMA_signal_3385, n3485}), .c ({new_AGEMA_signal_3661, n3624}) ) ;
    xnor_HPC2 U3506 ( .a ({new_AGEMA_signal_3945, n3392}), .b ({new_AGEMA_signal_3661, n3624}), .c ({state_out_s1[260], state_out_s0[260]}) ) ;
    xnor_HPC2 U3507 ( .a ({new_AGEMA_signal_3600, n3660}), .b ({new_AGEMA_signal_3654, n3656}), .c ({new_AGEMA_signal_3946, n3393}) ) ;
    xnor_HPC2 U3508 ( .a ({new_AGEMA_signal_3946, n3393}), .b ({new_AGEMA_signal_3661, n3624}), .c ({state_out_s1[299], state_out_s0[299]}) ) ;
    xnor_HPC2 U3509 ( .a ({new_AGEMA_signal_3336, n3395}), .b ({new_AGEMA_signal_3331, n3394}), .c ({new_AGEMA_signal_3662, n3846}) ) ;
    xnor_HPC2 U3510 ( .a ({new_AGEMA_signal_3645, n3637}), .b ({new_AGEMA_signal_3662, n3846}), .c ({new_AGEMA_signal_3947, n3397}) ) ;
    xor_HPC2 U3511 ( .a ({new_AGEMA_signal_3230, z0[10]}), .b ({state_in_s1[50], state_in_s0[50]}), .c ({new_AGEMA_signal_3386, n3398}) ) ;
    xnor_HPC2 U3512 ( .a ({new_AGEMA_signal_3386, n3398}), .b ({new_AGEMA_signal_3304, n3396}), .c ({new_AGEMA_signal_3663, n3843}) ) ;
    xnor_HPC2 U3513 ( .a ({new_AGEMA_signal_3947, n3397}), .b ({new_AGEMA_signal_3663, n3843}), .c ({state_out_s1[15], state_out_s0[15]}) ) ;
    xor_HPC2 U3514 ( .a ({new_AGEMA_signal_2991, z1[10]}), .b ({state_in_s1[306], state_in_s0[306]}), .c ({new_AGEMA_signal_3387, n3400}) ) ;
    xnor_HPC2 U3515 ( .a ({state_in_s1[114], state_in_s0[114]}), .b ({new_AGEMA_signal_3386, n3398}), .c ({new_AGEMA_signal_3664, n3399}) ) ;
    xnor_HPC2 U3516 ( .a ({new_AGEMA_signal_3387, n3400}), .b ({new_AGEMA_signal_3664, n3399}), .c ({new_AGEMA_signal_3948, n3884}) ) ;
    xnor_HPC2 U3517 ( .a ({new_AGEMA_signal_3918, n3412}), .b ({new_AGEMA_signal_3948, n3884}), .c ({new_AGEMA_signal_4246, n3403}) ) ;
    xor_HPC2 U3518 ( .a ({new_AGEMA_signal_3013, z1[32]}), .b ({state_in_s1[280], state_in_s0[280]}), .c ({new_AGEMA_signal_3388, n3402}) ) ;
    xor_HPC2 U3519 ( .a ({new_AGEMA_signal_3268, z0[32]}), .b ({state_in_s1[24], state_in_s0[24]}), .c ({new_AGEMA_signal_3389, n3604}) ) ;
    xnor_HPC2 U3520 ( .a ({state_in_s1[88], state_in_s0[88]}), .b ({new_AGEMA_signal_3389, n3604}), .c ({new_AGEMA_signal_3665, n3401}) ) ;
    xnor_HPC2 U3521 ( .a ({new_AGEMA_signal_3388, n3402}), .b ({new_AGEMA_signal_3665, n3401}), .c ({new_AGEMA_signal_3949, n3878}) ) ;
    xnor_HPC2 U3522 ( .a ({new_AGEMA_signal_4246, n3403}), .b ({new_AGEMA_signal_3949, n3878}), .c ({state_out_s1[91], state_out_s0[91]}) ) ;
    xor_HPC2 U3523 ( .a ({new_AGEMA_signal_3231, z0[13]}), .b ({state_in_s1[53], state_in_s0[53]}), .c ({new_AGEMA_signal_3390, n3413}) ) ;
    xnor_HPC2 U3524 ( .a ({new_AGEMA_signal_3390, n3413}), .b ({new_AGEMA_signal_3317, n3404}), .c ({new_AGEMA_signal_3666, n3887}) ) ;
    xor_HPC2 U3525 ( .a ({new_AGEMA_signal_3243, z0[22]}), .b ({state_in_s1[46], state_in_s0[46]}), .c ({new_AGEMA_signal_3391, n3546}) ) ;
    xnor_HPC2 U3526 ( .a ({new_AGEMA_signal_3391, n3546}), .b ({new_AGEMA_signal_3295, n3405}), .c ({new_AGEMA_signal_3667, n3806}) ) ;
    xnor_HPC2 U3527 ( .a ({new_AGEMA_signal_3666, n3887}), .b ({new_AGEMA_signal_3667, n3806}), .c ({new_AGEMA_signal_3950, n3408}) ) ;
    xnor_HPC2 U3528 ( .a ({new_AGEMA_signal_3332, n3407}), .b ({new_AGEMA_signal_3362, n3406}), .c ({new_AGEMA_signal_3668, n3803}) ) ;
    xnor_HPC2 U3529 ( .a ({new_AGEMA_signal_3950, n3408}), .b ({new_AGEMA_signal_3668, n3803}), .c ({state_out_s1[2], state_out_s0[2]}) ) ;
    xor_HPC2 U3530 ( .a ({new_AGEMA_signal_3019, z1[38]}), .b ({state_in_s1[286], state_in_s0[286]}), .c ({new_AGEMA_signal_3392, n3411}) ) ;
    xnor_HPC2 U3531 ( .a ({state_in_s1[94], state_in_s0[94]}), .b ({new_AGEMA_signal_3363, n3409}), .c ({new_AGEMA_signal_3669, n3410}) ) ;
    xnor_HPC2 U3532 ( .a ({new_AGEMA_signal_3392, n3411}), .b ({new_AGEMA_signal_3669, n3410}), .c ({new_AGEMA_signal_3951, n3607}) ) ;
    xnor_HPC2 U3533 ( .a ({new_AGEMA_signal_3918, n3412}), .b ({new_AGEMA_signal_3951, n3607}), .c ({new_AGEMA_signal_4248, n3416}) ) ;
    xor_HPC2 U3534 ( .a ({new_AGEMA_signal_2994, z1[13]}), .b ({state_in_s1[309], state_in_s0[309]}), .c ({new_AGEMA_signal_3393, n3415}) ) ;
    xnor_HPC2 U3535 ( .a ({state_in_s1[117], state_in_s0[117]}), .b ({new_AGEMA_signal_3390, n3413}), .c ({new_AGEMA_signal_3670, n3414}) ) ;
    xnor_HPC2 U3536 ( .a ({new_AGEMA_signal_3393, n3415}), .b ({new_AGEMA_signal_3670, n3414}), .c ({new_AGEMA_signal_3952, n3435}) ) ;
    xnor_HPC2 U3537 ( .a ({new_AGEMA_signal_4248, n3416}), .b ({new_AGEMA_signal_3952, n3435}), .c ({state_out_s1[94], state_out_s0[94]}) ) ;
    xnor_HPC2 U3538 ( .a ({new_AGEMA_signal_3909, n3433}), .b ({new_AGEMA_signal_3922, n3608}), .c ({new_AGEMA_signal_4249, n3417}) ) ;
    xnor_HPC2 U3539 ( .a ({new_AGEMA_signal_4249, n3417}), .b ({new_AGEMA_signal_3952, n3435}), .c ({state_out_s1[104], state_out_s0[104]}) ) ;
    xor_HPC2 U3540 ( .a ({new_AGEMA_signal_3257, z0[27]}), .b ({state_in_s1[35], state_in_s0[35]}), .c ({new_AGEMA_signal_3394, n3427}) ) ;
    xnor_HPC2 U3541 ( .a ({state_in_s1[227], state_in_s0[227]}), .b ({new_AGEMA_signal_3130, z4[27]}), .c ({new_AGEMA_signal_3395, n3423}) ) ;
    xnor_HPC2 U3542 ( .a ({new_AGEMA_signal_3394, n3427}), .b ({new_AGEMA_signal_3395, n3423}), .c ({new_AGEMA_signal_3671, n3856}) ) ;
    xor_HPC2 U3543 ( .a ({new_AGEMA_signal_3262, z0[36]}), .b ({state_in_s1[28], state_in_s0[28]}), .c ({new_AGEMA_signal_3396, n3444}) ) ;
    xnor_HPC2 U3544 ( .a ({new_AGEMA_signal_3396, n3444}), .b ({new_AGEMA_signal_3327, n3418}), .c ({new_AGEMA_signal_3672, n3787}) ) ;
    xnor_HPC2 U3545 ( .a ({new_AGEMA_signal_3671, n3856}), .b ({new_AGEMA_signal_3672, n3787}), .c ({new_AGEMA_signal_3953, n3421}) ) ;
    xnor_HPC2 U3546 ( .a ({new_AGEMA_signal_3369, n3420}), .b ({new_AGEMA_signal_3298, n3419}), .c ({new_AGEMA_signal_3673, n3774}) ) ;
    xnor_HPC2 U3547 ( .a ({new_AGEMA_signal_3953, n3421}), .b ({new_AGEMA_signal_3673, n3774}), .c ({state_out_s1[48], state_out_s0[48]}) ) ;
    xnor_HPC2 U3548 ( .a ({new_AGEMA_signal_3599, n3454}), .b ({new_AGEMA_signal_3615, n3422}), .c ({new_AGEMA_signal_3954, n3424}) ) ;
    xnor_HPC2 U3549 ( .a ({state_in_s1[291], state_in_s0[291]}), .b ({new_AGEMA_signal_3395, n3423}), .c ({new_AGEMA_signal_3674, n3725}) ) ;
    xnor_HPC2 U3550 ( .a ({new_AGEMA_signal_3954, n3424}), .b ({new_AGEMA_signal_3674, n3725}), .c ({state_out_s1[291], state_out_s0[291]}) ) ;
    xor_HPC2 U3551 ( .a ({new_AGEMA_signal_3030, z1[49]}), .b ({state_in_s1[265], state_in_s0[265]}), .c ({new_AGEMA_signal_3397, n3426}) ) ;
    xor_HPC2 U3552 ( .a ({new_AGEMA_signal_3237, z0[49]}), .b ({state_in_s1[9], state_in_s0[9]}), .c ({new_AGEMA_signal_3398, n3653}) ) ;
    xnor_HPC2 U3553 ( .a ({state_in_s1[73], state_in_s0[73]}), .b ({new_AGEMA_signal_3398, n3653}), .c ({new_AGEMA_signal_3675, n3425}) ) ;
    xnor_HPC2 U3554 ( .a ({new_AGEMA_signal_3397, n3426}), .b ({new_AGEMA_signal_3675, n3425}), .c ({new_AGEMA_signal_3955, n3883}) ) ;
    xor_HPC2 U3555 ( .a ({new_AGEMA_signal_3008, z1[27]}), .b ({state_in_s1[291], state_in_s0[291]}), .c ({new_AGEMA_signal_3399, n3429}) ) ;
    xnor_HPC2 U3556 ( .a ({state_in_s1[99], state_in_s0[99]}), .b ({new_AGEMA_signal_3394, n3427}), .c ({new_AGEMA_signal_3676, n3428}) ) ;
    xnor_HPC2 U3557 ( .a ({new_AGEMA_signal_3399, n3429}), .b ({new_AGEMA_signal_3676, n3428}), .c ({new_AGEMA_signal_3956, n3744}) ) ;
    xnor_HPC2 U3558 ( .a ({new_AGEMA_signal_3955, n3883}), .b ({new_AGEMA_signal_3956, n3744}), .c ({new_AGEMA_signal_4252, n3432}) ) ;
    xor_HPC2 U3559 ( .a ({new_AGEMA_signal_3232, z0[52]}), .b ({state_in_s1[12], state_in_s0[12]}), .c ({new_AGEMA_signal_3400, n3912}) ) ;
    xor_HPC2 U3560 ( .a ({new_AGEMA_signal_3033, z1[52]}), .b ({new_AGEMA_signal_3400, n3912}), .c ({new_AGEMA_signal_3677, n3431}) ) ;
    xnor_HPC2 U3562 ( .a ({new_AGEMA_signal_3677, n3431}), .b ({new_AGEMA_signal_2675, n3430}), .c ({new_AGEMA_signal_3957, n3436}) ) ;
    xnor_HPC2 U3563 ( .a ({new_AGEMA_signal_4252, n3432}), .b ({new_AGEMA_signal_3957, n3436}), .c ({state_out_s1[76], state_out_s0[76]}) ) ;
    xnor_HPC2 U3564 ( .a ({new_AGEMA_signal_3909, n3433}), .b ({new_AGEMA_signal_3933, n3745}), .c ({new_AGEMA_signal_4253, n3434}) ) ;
    xnor_HPC2 U3565 ( .a ({new_AGEMA_signal_4253, n3434}), .b ({new_AGEMA_signal_3957, n3436}), .c ({state_out_s1[79], state_out_s0[79]}) ) ;
    xnor_HPC2 U3566 ( .a ({new_AGEMA_signal_3948, n3884}), .b ({new_AGEMA_signal_3952, n3435}), .c ({new_AGEMA_signal_4254, n3437}) ) ;
    xnor_HPC2 U3567 ( .a ({new_AGEMA_signal_4254, n3437}), .b ({new_AGEMA_signal_3957, n3436}), .c ({state_out_s1[117], state_out_s0[117]}) ) ;
    xor_HPC2 U3568 ( .a ({new_AGEMA_signal_3227, z0[11]}), .b ({state_in_s1[51], state_in_s0[51]}), .c ({new_AGEMA_signal_3401, n3448}) ) ;
    xnor_HPC2 U3569 ( .a ({new_AGEMA_signal_3401, n3448}), .b ({new_AGEMA_signal_3307, n3438}), .c ({new_AGEMA_signal_3678, n3704}) ) ;
    xnor_HPC2 U3570 ( .a ({new_AGEMA_signal_3360, n3440}), .b ({new_AGEMA_signal_3315, n3439}), .c ({new_AGEMA_signal_3679, n3671}) ) ;
    xnor_HPC2 U3571 ( .a ({new_AGEMA_signal_3678, n3704}), .b ({new_AGEMA_signal_3679, n3671}), .c ({new_AGEMA_signal_3958, n3443}) ) ;
    xnor_HPC2 U3572 ( .a ({new_AGEMA_signal_3341, n3442}), .b ({new_AGEMA_signal_3297, n3441}), .c ({new_AGEMA_signal_3680, n3667}) ) ;
    xnor_HPC2 U3573 ( .a ({new_AGEMA_signal_3958, n3443}), .b ({new_AGEMA_signal_3680, n3667}), .c ({state_out_s1[0], state_out_s0[0]}) ) ;
    xor_HPC2 U3574 ( .a ({new_AGEMA_signal_3017, z1[36]}), .b ({state_in_s1[284], state_in_s0[284]}), .c ({new_AGEMA_signal_3402, n3446}) ) ;
    xnor_HPC2 U3575 ( .a ({state_in_s1[92], state_in_s0[92]}), .b ({new_AGEMA_signal_3396, n3444}), .c ({new_AGEMA_signal_3681, n3445}) ) ;
    xnor_HPC2 U3576 ( .a ({new_AGEMA_signal_3402, n3446}), .b ({new_AGEMA_signal_3681, n3445}), .c ({new_AGEMA_signal_3959, n3541}) ) ;
    xnor_HPC2 U3577 ( .a ({new_AGEMA_signal_3908, n3447}), .b ({new_AGEMA_signal_3959, n3541}), .c ({new_AGEMA_signal_4256, n3451}) ) ;
    xor_HPC2 U3578 ( .a ({new_AGEMA_signal_2992, z1[11]}), .b ({new_AGEMA_signal_3401, n3448}), .c ({new_AGEMA_signal_3682, n3450}) ) ;
    xnor_HPC2 U3580 ( .a ({new_AGEMA_signal_3682, n3450}), .b ({new_AGEMA_signal_2677, n3449}), .c ({new_AGEMA_signal_3960, n3472}) ) ;
    xnor_HPC2 U3581 ( .a ({new_AGEMA_signal_4256, n3451}), .b ({new_AGEMA_signal_3960, n3472}), .c ({state_out_s1[92], state_out_s0[92]}) ) ;
    xnor_HPC2 U3582 ( .a ({new_AGEMA_signal_3932, n3751}), .b ({new_AGEMA_signal_3936, n3468}), .c ({new_AGEMA_signal_4257, n3452}) ) ;
    xnor_HPC2 U3583 ( .a ({new_AGEMA_signal_4257, n3452}), .b ({new_AGEMA_signal_3960, n3472}), .c ({state_out_s1[115], state_out_s0[115]}) ) ;
    xnor_HPC2 U3584 ( .a ({new_AGEMA_signal_3599, n3454}), .b ({new_AGEMA_signal_3628, n3453}), .c ({new_AGEMA_signal_3961, n3455}) ) ;
    xnor_HPC2 U3585 ( .a ({state_in_s1[197], state_in_s0[197]}), .b ({new_AGEMA_signal_3168, z4[61]}), .c ({new_AGEMA_signal_3403, n3680}) ) ;
    xnor_HPC2 U3586 ( .a ({state_in_s1[261], state_in_s0[261]}), .b ({new_AGEMA_signal_3403, n3680}), .c ({new_AGEMA_signal_3683, n3459}) ) ;
    xnor_HPC2 U3587 ( .a ({new_AGEMA_signal_3961, n3455}), .b ({new_AGEMA_signal_3683, n3459}), .c ({state_out_s1[261], state_out_s0[261]}) ) ;
    xnor_HPC2 U3588 ( .a ({new_AGEMA_signal_3606, n3457}), .b ({new_AGEMA_signal_3629, n3456}), .c ({new_AGEMA_signal_3962, n3458}) ) ;
    xnor_HPC2 U3589 ( .a ({new_AGEMA_signal_3962, n3458}), .b ({new_AGEMA_signal_3683, n3459}), .c ({state_out_s1[270], state_out_s0[270]}) ) ;
    xnor_HPC2 U3590 ( .a ({new_AGEMA_signal_3605, n3729}), .b ({new_AGEMA_signal_3674, n3725}), .c ({new_AGEMA_signal_3963, n3460}) ) ;
    xnor_HPC2 U3591 ( .a ({new_AGEMA_signal_3963, n3460}), .b ({new_AGEMA_signal_3683, n3459}), .c ({state_out_s1[300], state_out_s0[300]}) ) ;
    xnor_HPC2 U3592 ( .a ({new_AGEMA_signal_3912, n3464}), .b ({new_AGEMA_signal_3926, n3617}), .c ({new_AGEMA_signal_4261, n3463}) ) ;
    xor_HPC2 U3593 ( .a ({new_AGEMA_signal_2995, z1[14]}), .b ({state_in_s1[310], state_in_s0[310]}), .c ({new_AGEMA_signal_3404, n3462}) ) ;
    xor_HPC2 U3594 ( .a ({new_AGEMA_signal_3228, z0[14]}), .b ({state_in_s1[54], state_in_s0[54]}), .c ({new_AGEMA_signal_3405, n3599}) ) ;
    xnor_HPC2 U3595 ( .a ({state_in_s1[118], state_in_s0[118]}), .b ({new_AGEMA_signal_3405, n3599}), .c ({new_AGEMA_signal_3684, n3461}) ) ;
    xnor_HPC2 U3596 ( .a ({new_AGEMA_signal_3404, n3462}), .b ({new_AGEMA_signal_3684, n3461}), .c ({new_AGEMA_signal_3964, n3530}) ) ;
    xnor_HPC2 U3597 ( .a ({new_AGEMA_signal_4261, n3463}), .b ({new_AGEMA_signal_3964, n3530}), .c ({state_out_s1[105], state_out_s0[105]}) ) ;
    xnor_HPC2 U3598 ( .a ({new_AGEMA_signal_3912, n3464}), .b ({new_AGEMA_signal_3941, n3762}), .c ({new_AGEMA_signal_4262, n3467}) ) ;
    xor_HPC2 U3599 ( .a ({new_AGEMA_signal_3034, z1[53]}), .b ({state_in_s1[269], state_in_s0[269]}), .c ({new_AGEMA_signal_3406, n3466}) ) ;
    xor_HPC2 U3600 ( .a ({new_AGEMA_signal_3229, z0[53]}), .b ({state_in_s1[13], state_in_s0[13]}), .c ({new_AGEMA_signal_3407, n3567}) ) ;
    xnor_HPC2 U3601 ( .a ({state_in_s1[77], state_in_s0[77]}), .b ({new_AGEMA_signal_3407, n3567}), .c ({new_AGEMA_signal_3685, n3465}) ) ;
    xnor_HPC2 U3602 ( .a ({new_AGEMA_signal_3406, n3466}), .b ({new_AGEMA_signal_3685, n3465}), .c ({new_AGEMA_signal_3965, n3473}) ) ;
    xnor_HPC2 U3603 ( .a ({new_AGEMA_signal_4262, n3467}), .b ({new_AGEMA_signal_3965, n3473}), .c ({state_out_s1[64], state_out_s0[64]}) ) ;
    xnor_HPC2 U3604 ( .a ({new_AGEMA_signal_3936, n3468}), .b ({new_AGEMA_signal_3965, n3473}), .c ({new_AGEMA_signal_4263, n3471}) ) ;
    xor_HPC2 U3605 ( .a ({new_AGEMA_signal_3255, z0[28]}), .b ({state_in_s1[36], state_in_s0[36]}), .c ({new_AGEMA_signal_3408, n3475}) ) ;
    xor_HPC2 U3606 ( .a ({new_AGEMA_signal_3009, z1[28]}), .b ({new_AGEMA_signal_3408, n3475}), .c ({new_AGEMA_signal_3686, n3470}) ) ;
    xnor_HPC2 U3608 ( .a ({new_AGEMA_signal_3686, n3470}), .b ({new_AGEMA_signal_2679, n3469}), .c ({new_AGEMA_signal_3966, n3809}) ) ;
    xnor_HPC2 U3609 ( .a ({new_AGEMA_signal_4263, n3471}), .b ({new_AGEMA_signal_3966, n3809}), .c ({state_out_s1[77], state_out_s0[77]}) ) ;
    xnor_HPC2 U3610 ( .a ({new_AGEMA_signal_3960, n3472}), .b ({new_AGEMA_signal_3964, n3530}), .c ({new_AGEMA_signal_4264, n3474}) ) ;
    xnor_HPC2 U3611 ( .a ({new_AGEMA_signal_4264, n3474}), .b ({new_AGEMA_signal_3965, n3473}), .c ({state_out_s1[118], state_out_s0[118]}) ) ;
    xnor_HPC2 U3612 ( .a ({new_AGEMA_signal_3644, n3705}), .b ({new_AGEMA_signal_3680, n3667}), .c ({new_AGEMA_signal_3967, n3476}) ) ;
    xnor_HPC2 U3613 ( .a ({state_in_s1[228], state_in_s0[228]}), .b ({new_AGEMA_signal_3131, z4[28]}), .c ({new_AGEMA_signal_3409, n3482}) ) ;
    xnor_HPC2 U3614 ( .a ({new_AGEMA_signal_3408, n3475}), .b ({new_AGEMA_signal_3409, n3482}), .c ({new_AGEMA_signal_3687, n3636}) ) ;
    xnor_HPC2 U3615 ( .a ({new_AGEMA_signal_3967, n3476}), .b ({new_AGEMA_signal_3687, n3636}), .c ({state_out_s1[36], state_out_s0[36]}) ) ;
    xor_HPC2 U3616 ( .a ({new_AGEMA_signal_3266, z0[37]}), .b ({state_in_s1[29], state_in_s0[29]}), .c ({new_AGEMA_signal_3410, n3499}) ) ;
    xnor_HPC2 U3617 ( .a ({new_AGEMA_signal_3410, n3499}), .b ({new_AGEMA_signal_3328, n3477}), .c ({new_AGEMA_signal_3688, n3863}) ) ;
    xnor_HPC2 U3618 ( .a ({new_AGEMA_signal_3687, n3636}), .b ({new_AGEMA_signal_3688, n3863}), .c ({new_AGEMA_signal_3968, n3480}) ) ;
    xnor_HPC2 U3619 ( .a ({new_AGEMA_signal_3378, n3479}), .b ({new_AGEMA_signal_3301, n3478}), .c ({new_AGEMA_signal_3689, n3860}) ) ;
    xnor_HPC2 U3620 ( .a ({new_AGEMA_signal_3968, n3480}), .b ({new_AGEMA_signal_3689, n3860}), .c ({state_out_s1[49], state_out_s0[49]}) ) ;
    xnor_HPC2 U3621 ( .a ({new_AGEMA_signal_3604, n3508}), .b ({new_AGEMA_signal_3616, n3481}), .c ({new_AGEMA_signal_3969, n3483}) ) ;
    xnor_HPC2 U3622 ( .a ({state_in_s1[292], state_in_s0[292]}), .b ({new_AGEMA_signal_3409, n3482}), .c ({new_AGEMA_signal_3690, n3831}) ) ;
    xnor_HPC2 U3623 ( .a ({new_AGEMA_signal_3969, n3483}), .b ({new_AGEMA_signal_3690, n3831}), .c ({state_out_s1[292], state_out_s0[292]}) ) ;
    xor_HPC2 U3624 ( .a ({new_AGEMA_signal_3261, z0[24]}), .b ({state_in_s1[32], state_in_s0[32]}), .c ({new_AGEMA_signal_3411, n3591}) ) ;
    xnor_HPC2 U3625 ( .a ({new_AGEMA_signal_3411, n3591}), .b ({new_AGEMA_signal_3358, n3484}), .c ({new_AGEMA_signal_3691, n3918}) ) ;
    xnor_HPC2 U3626 ( .a ({new_AGEMA_signal_3347, n3486}), .b ({new_AGEMA_signal_3385, n3485}), .c ({new_AGEMA_signal_3692, n3826}) ) ;
    xnor_HPC2 U3627 ( .a ({new_AGEMA_signal_3691, n3918}), .b ({new_AGEMA_signal_3692, n3826}), .c ({new_AGEMA_signal_3970, n3488}) ) ;
    xor_HPC2 U3628 ( .a ({new_AGEMA_signal_3224, z0[15]}), .b ({state_in_s1[55], state_in_s0[55]}), .c ({new_AGEMA_signal_3412, n3489}) ) ;
    xnor_HPC2 U3629 ( .a ({new_AGEMA_signal_3412, n3489}), .b ({new_AGEMA_signal_3296, n3487}), .c ({new_AGEMA_signal_3693, n3823}) ) ;
    xnor_HPC2 U3630 ( .a ({new_AGEMA_signal_3970, n3488}), .b ({new_AGEMA_signal_3693, n3823}), .c ({state_out_s1[4], state_out_s0[4]}) ) ;
    xnor_HPC2 U3631 ( .a ({new_AGEMA_signal_3917, n3515}), .b ({new_AGEMA_signal_3920, n3648}), .c ({new_AGEMA_signal_4269, n3492}) ) ;
    xor_HPC2 U3632 ( .a ({new_AGEMA_signal_2996, z1[15]}), .b ({state_in_s1[311], state_in_s0[311]}), .c ({new_AGEMA_signal_3413, n3491}) ) ;
    xnor_HPC2 U3633 ( .a ({state_in_s1[119], state_in_s0[119]}), .b ({new_AGEMA_signal_3412, n3489}), .c ({new_AGEMA_signal_3694, n3490}) ) ;
    xnor_HPC2 U3634 ( .a ({new_AGEMA_signal_3413, n3491}), .b ({new_AGEMA_signal_3694, n3490}), .c ({new_AGEMA_signal_3971, n3554}) ) ;
    xnor_HPC2 U3635 ( .a ({new_AGEMA_signal_4269, n3492}), .b ({new_AGEMA_signal_3971, n3554}), .c ({state_out_s1[106], state_out_s0[106]}) ) ;
    xor_HPC2 U3636 ( .a ({new_AGEMA_signal_3225, z0[12]}), .b ({state_in_s1[52], state_in_s0[52]}), .c ({new_AGEMA_signal_3414, n3503}) ) ;
    xnor_HPC2 U3637 ( .a ({new_AGEMA_signal_3414, n3503}), .b ({new_AGEMA_signal_3312, n3493}), .c ({new_AGEMA_signal_3695, n3799}) ) ;
    xnor_HPC2 U3638 ( .a ({new_AGEMA_signal_3352, n3495}), .b ({new_AGEMA_signal_3330, n3494}), .c ({new_AGEMA_signal_3696, n3712}) ) ;
    xnor_HPC2 U3639 ( .a ({new_AGEMA_signal_3695, n3799}), .b ({new_AGEMA_signal_3696, n3712}), .c ({new_AGEMA_signal_3972, n3498}) ) ;
    xnor_HPC2 U3640 ( .a ({new_AGEMA_signal_3348, n3497}), .b ({new_AGEMA_signal_3344, n3496}), .c ({new_AGEMA_signal_3697, n3708}) ) ;
    xnor_HPC2 U3641 ( .a ({new_AGEMA_signal_3972, n3498}), .b ({new_AGEMA_signal_3697, n3708}), .c ({state_out_s1[1], state_out_s0[1]}) ) ;
    xor_HPC2 U3642 ( .a ({new_AGEMA_signal_3018, z1[37]}), .b ({state_in_s1[285], state_in_s0[285]}), .c ({new_AGEMA_signal_3415, n3501}) ) ;
    xnor_HPC2 U3643 ( .a ({state_in_s1[93], state_in_s0[93]}), .b ({new_AGEMA_signal_3410, n3499}), .c ({new_AGEMA_signal_3698, n3500}) ) ;
    xnor_HPC2 U3644 ( .a ({new_AGEMA_signal_3415, n3501}), .b ({new_AGEMA_signal_3698, n3500}), .c ({new_AGEMA_signal_3973, n3571}) ) ;
    xnor_HPC2 U3645 ( .a ({new_AGEMA_signal_3911, n3502}), .b ({new_AGEMA_signal_3973, n3571}), .c ({new_AGEMA_signal_4271, n3506}) ) ;
    xor_HPC2 U3646 ( .a ({new_AGEMA_signal_2993, z1[12]}), .b ({state_in_s1[308], state_in_s0[308]}), .c ({new_AGEMA_signal_3416, n3505}) ) ;
    xnor_HPC2 U3647 ( .a ({state_in_s1[116], state_in_s0[116]}), .b ({new_AGEMA_signal_3414, n3503}), .c ({new_AGEMA_signal_3699, n3504}) ) ;
    xnor_HPC2 U3648 ( .a ({new_AGEMA_signal_3416, n3505}), .b ({new_AGEMA_signal_3699, n3504}), .c ({new_AGEMA_signal_3974, n3523}) ) ;
    xnor_HPC2 U3649 ( .a ({new_AGEMA_signal_4271, n3506}), .b ({new_AGEMA_signal_3974, n3523}), .c ({state_out_s1[93], state_out_s0[93]}) ) ;
    xnor_HPC2 U3650 ( .a ({new_AGEMA_signal_3940, n3767}), .b ({new_AGEMA_signal_3944, n3519}), .c ({new_AGEMA_signal_4272, n3507}) ) ;
    xnor_HPC2 U3651 ( .a ({new_AGEMA_signal_4272, n3507}), .b ({new_AGEMA_signal_3974, n3523}), .c ({state_out_s1[116], state_out_s0[116]}) ) ;
    xnor_HPC2 U3652 ( .a ({new_AGEMA_signal_3604, n3508}), .b ({new_AGEMA_signal_3610, n3686}), .c ({new_AGEMA_signal_3975, n3509}) ) ;
    xnor_HPC2 U3653 ( .a ({state_in_s1[198], state_in_s0[198]}), .b ({new_AGEMA_signal_3169, z4[62]}), .c ({new_AGEMA_signal_3417, n3565}) ) ;
    xnor_HPC2 U3654 ( .a ({state_in_s1[262], state_in_s0[262]}), .b ({new_AGEMA_signal_3417, n3565}), .c ({new_AGEMA_signal_3700, n3513}) ) ;
    xnor_HPC2 U3655 ( .a ({new_AGEMA_signal_3975, n3509}), .b ({new_AGEMA_signal_3700, n3513}), .c ({state_out_s1[262], state_out_s0[262]}) ) ;
    xnor_HPC2 U3656 ( .a ({new_AGEMA_signal_3611, n3511}), .b ({new_AGEMA_signal_3621, n3510}), .c ({new_AGEMA_signal_3976, n3512}) ) ;
    xnor_HPC2 U3657 ( .a ({new_AGEMA_signal_3976, n3512}), .b ({new_AGEMA_signal_3700, n3513}), .c ({state_out_s1[271], state_out_s0[271]}) ) ;
    xnor_HPC2 U3658 ( .a ({new_AGEMA_signal_3620, n3835}), .b ({new_AGEMA_signal_3690, n3831}), .c ({new_AGEMA_signal_3977, n3514}) ) ;
    xnor_HPC2 U3659 ( .a ({new_AGEMA_signal_3977, n3514}), .b ({new_AGEMA_signal_3700, n3513}), .c ({state_out_s1[301], state_out_s0[301]}) ) ;
    xnor_HPC2 U3660 ( .a ({new_AGEMA_signal_3917, n3515}), .b ({new_AGEMA_signal_3949, n3878}), .c ({new_AGEMA_signal_4276, n3518}) ) ;
    xor_HPC2 U3661 ( .a ({new_AGEMA_signal_3035, z1[54]}), .b ({state_in_s1[270], state_in_s0[270]}), .c ({new_AGEMA_signal_3418, n3517}) ) ;
    xor_HPC2 U3662 ( .a ({new_AGEMA_signal_3226, z0[54]}), .b ({state_in_s1[14], state_in_s0[14]}), .c ({new_AGEMA_signal_3419, n3583}) ) ;
    xnor_HPC2 U3663 ( .a ({state_in_s1[78], state_in_s0[78]}), .b ({new_AGEMA_signal_3419, n3583}), .c ({new_AGEMA_signal_3701, n3516}) ) ;
    xnor_HPC2 U3664 ( .a ({new_AGEMA_signal_3418, n3517}), .b ({new_AGEMA_signal_3701, n3516}), .c ({new_AGEMA_signal_3978, n3524}) ) ;
    xnor_HPC2 U3665 ( .a ({new_AGEMA_signal_4276, n3518}), .b ({new_AGEMA_signal_3978, n3524}), .c ({state_out_s1[65], state_out_s0[65]}) ) ;
    xnor_HPC2 U3666 ( .a ({new_AGEMA_signal_3944, n3519}), .b ({new_AGEMA_signal_3978, n3524}), .c ({new_AGEMA_signal_4277, n3522}) ) ;
    xor_HPC2 U3667 ( .a ({new_AGEMA_signal_3259, z0[29]}), .b ({state_in_s1[37], state_in_s0[37]}), .c ({new_AGEMA_signal_3420, n3535}) ) ;
    xor_HPC2 U3668 ( .a ({new_AGEMA_signal_3010, z1[29]}), .b ({new_AGEMA_signal_3420, n3535}), .c ({new_AGEMA_signal_3702, n3521}) ) ;
    xnor_HPC2 U3670 ( .a ({new_AGEMA_signal_3702, n3521}), .b ({new_AGEMA_signal_2681, n3520}), .c ({new_AGEMA_signal_3979, n3897}) ) ;
    xnor_HPC2 U3671 ( .a ({new_AGEMA_signal_4277, n3522}), .b ({new_AGEMA_signal_3979, n3897}), .c ({state_out_s1[78], state_out_s0[78]}) ) ;
    xnor_HPC2 U3672 ( .a ({new_AGEMA_signal_3971, n3554}), .b ({new_AGEMA_signal_3974, n3523}), .c ({new_AGEMA_signal_4278, n3525}) ) ;
    xnor_HPC2 U3673 ( .a ({new_AGEMA_signal_4278, n3525}), .b ({new_AGEMA_signal_3978, n3524}), .c ({state_out_s1[119], state_out_s0[119]}) ) ;
    xor_HPC2 U3674 ( .a ({new_AGEMA_signal_3222, z0[39]}), .b ({state_in_s1[31], state_in_s0[31]}), .c ({new_AGEMA_signal_3421, n3531}) ) ;
    xnor_HPC2 U3675 ( .a ({new_AGEMA_signal_3421, n3531}), .b ({new_AGEMA_signal_3320, n3526}), .c ({new_AGEMA_signal_3703, n3802}) ) ;
    xnor_HPC2 U3676 ( .a ({new_AGEMA_signal_3679, n3671}), .b ({new_AGEMA_signal_3703, n3802}), .c ({new_AGEMA_signal_3980, n3529}) ) ;
    xnor_HPC2 U3677 ( .a ({new_AGEMA_signal_3383, n3528}), .b ({new_AGEMA_signal_3366, n3527}), .c ({new_AGEMA_signal_3704, n3798}) ) ;
    xnor_HPC2 U3678 ( .a ({new_AGEMA_signal_3980, n3529}), .b ({new_AGEMA_signal_3704, n3798}), .c ({state_out_s1[44], state_out_s0[44]}) ) ;
    xnor_HPC2 U3679 ( .a ({new_AGEMA_signal_3959, n3541}), .b ({new_AGEMA_signal_3964, n3530}), .c ({new_AGEMA_signal_4280, n3534}) ) ;
    xor_HPC2 U3680 ( .a ({new_AGEMA_signal_3020, z1[39]}), .b ({state_in_s1[287], state_in_s0[287]}), .c ({new_AGEMA_signal_3422, n3533}) ) ;
    xnor_HPC2 U3681 ( .a ({state_in_s1[95], state_in_s0[95]}), .b ({new_AGEMA_signal_3421, n3531}), .c ({new_AGEMA_signal_3705, n3532}) ) ;
    xnor_HPC2 U3682 ( .a ({new_AGEMA_signal_3422, n3533}), .b ({new_AGEMA_signal_3705, n3532}), .c ({new_AGEMA_signal_3981, n3644}) ) ;
    xnor_HPC2 U3683 ( .a ({new_AGEMA_signal_4280, n3534}), .b ({new_AGEMA_signal_3981, n3644}), .c ({state_out_s1[95], state_out_s0[95]}) ) ;
    xnor_HPC2 U3684 ( .a ({new_AGEMA_signal_3697, n3708}), .b ({new_AGEMA_signal_3704, n3798}), .c ({new_AGEMA_signal_3982, n3536}) ) ;
    xnor_HPC2 U3685 ( .a ({state_in_s1[229], state_in_s0[229]}), .b ({new_AGEMA_signal_3132, z4[29]}), .c ({new_AGEMA_signal_3423, n3539}) ) ;
    xnor_HPC2 U3686 ( .a ({new_AGEMA_signal_3420, n3535}), .b ({new_AGEMA_signal_3423, n3539}), .c ({new_AGEMA_signal_3706, n3670}) ) ;
    xnor_HPC2 U3687 ( .a ({new_AGEMA_signal_3982, n3536}), .b ({new_AGEMA_signal_3706, n3670}), .c ({state_out_s1[37], state_out_s0[37]}) ) ;
    xnor_HPC2 U3688 ( .a ({new_AGEMA_signal_3643, n3709}), .b ({new_AGEMA_signal_3663, n3843}), .c ({new_AGEMA_signal_3983, n3537}) ) ;
    xnor_HPC2 U3689 ( .a ({new_AGEMA_signal_3983, n3537}), .b ({new_AGEMA_signal_3706, n3670}), .c ({state_out_s1[50], state_out_s0[50]}) ) ;
    xnor_HPC2 U3690 ( .a ({new_AGEMA_signal_3609, n3561}), .b ({new_AGEMA_signal_3617, n3538}), .c ({new_AGEMA_signal_3984, n3540}) ) ;
    xnor_HPC2 U3691 ( .a ({state_in_s1[293], state_in_s0[293]}), .b ({new_AGEMA_signal_3423, n3539}), .c ({new_AGEMA_signal_3707, n3921}) ) ;
    xnor_HPC2 U3692 ( .a ({new_AGEMA_signal_3984, n3540}), .b ({new_AGEMA_signal_3707, n3921}), .c ({state_out_s1[293], state_out_s0[293]}) ) ;
    xnor_HPC2 U3693 ( .a ({new_AGEMA_signal_3907, n3542}), .b ({new_AGEMA_signal_3959, n3541}), .c ({new_AGEMA_signal_4284, n3545}) ) ;
    xor_HPC2 U3694 ( .a ({new_AGEMA_signal_3042, z1[61]}), .b ({state_in_s1[261], state_in_s0[261]}), .c ({new_AGEMA_signal_3424, n3544}) ) ;
    xor_HPC2 U3695 ( .a ({new_AGEMA_signal_3223, z0[61]}), .b ({state_in_s1[5], state_in_s0[5]}), .c ({new_AGEMA_signal_3425, n3681}) ) ;
    xnor_HPC2 U3696 ( .a ({state_in_s1[69], state_in_s0[69]}), .b ({new_AGEMA_signal_3425, n3681}), .c ({new_AGEMA_signal_3708, n3543}) ) ;
    xnor_HPC2 U3697 ( .a ({new_AGEMA_signal_3424, n3544}), .b ({new_AGEMA_signal_3708, n3543}), .c ({new_AGEMA_signal_3985, n3643}) ) ;
    xnor_HPC2 U3698 ( .a ({new_AGEMA_signal_4284, n3545}), .b ({new_AGEMA_signal_3985, n3643}), .c ({state_out_s1[69], state_out_s0[69]}) ) ;
    xnor_HPC2 U3699 ( .a ({new_AGEMA_signal_3921, n3697}), .b ({new_AGEMA_signal_3985, n3643}), .c ({new_AGEMA_signal_4285, n3549}) ) ;
    xor_HPC2 U3700 ( .a ({new_AGEMA_signal_3003, z1[22]}), .b ({new_AGEMA_signal_3391, n3546}), .c ({new_AGEMA_signal_3709, n3548}) ) ;
    xnor_HPC2 U3702 ( .a ({new_AGEMA_signal_3709, n3548}), .b ({new_AGEMA_signal_2683, n3547}), .c ({new_AGEMA_signal_3986, n3702}) ) ;
    xnor_HPC2 U3703 ( .a ({new_AGEMA_signal_4285, n3549}), .b ({new_AGEMA_signal_3986, n3702}), .c ({state_out_s1[110], state_out_s0[110]}) ) ;
    xor_HPC2 U3704 ( .a ({new_AGEMA_signal_3220, z0[40]}), .b ({state_in_s1[16], state_in_s0[16]}), .c ({new_AGEMA_signal_3426, n3555}) ) ;
    xnor_HPC2 U3705 ( .a ({new_AGEMA_signal_3426, n3555}), .b ({new_AGEMA_signal_3322, n3550}), .c ({new_AGEMA_signal_3710, n3891}) ) ;
    xnor_HPC2 U3706 ( .a ({new_AGEMA_signal_3695, n3799}), .b ({new_AGEMA_signal_3710, n3891}), .c ({new_AGEMA_signal_3987, n3553}) ) ;
    xnor_HPC2 U3707 ( .a ({new_AGEMA_signal_3380, n3552}), .b ({new_AGEMA_signal_3343, n3551}), .c ({new_AGEMA_signal_3711, n3805}) ) ;
    xnor_HPC2 U3708 ( .a ({new_AGEMA_signal_3987, n3553}), .b ({new_AGEMA_signal_3711, n3805}), .c ({state_out_s1[52], state_out_s0[52]}) ) ;
    xnor_HPC2 U3709 ( .a ({new_AGEMA_signal_3971, n3554}), .b ({new_AGEMA_signal_3973, n3571}), .c ({new_AGEMA_signal_4287, n3558}) ) ;
    xor_HPC2 U3710 ( .a ({new_AGEMA_signal_3021, z1[40]}), .b ({state_in_s1[272], state_in_s0[272]}), .c ({new_AGEMA_signal_3427, n3557}) ) ;
    xnor_HPC2 U3711 ( .a ({state_in_s1[80], state_in_s0[80]}), .b ({new_AGEMA_signal_3426, n3555}), .c ({new_AGEMA_signal_3712, n3556}) ) ;
    xnor_HPC2 U3712 ( .a ({new_AGEMA_signal_3427, n3557}), .b ({new_AGEMA_signal_3712, n3556}), .c ({new_AGEMA_signal_3988, n3678}) ) ;
    xnor_HPC2 U3713 ( .a ({new_AGEMA_signal_4287, n3558}), .b ({new_AGEMA_signal_3988, n3678}), .c ({state_out_s1[80], state_out_s0[80]}) ) ;
    xnor_HPC2 U3714 ( .a ({new_AGEMA_signal_3587, n3657}), .b ({new_AGEMA_signal_3613, n3559}), .c ({new_AGEMA_signal_3989, n3560}) ) ;
    xnor_HPC2 U3715 ( .a ({state_in_s1[199], state_in_s0[199]}), .b ({new_AGEMA_signal_3170, z4[63]}), .c ({new_AGEMA_signal_3428, n3584}) ) ;
    xnor_HPC2 U3716 ( .a ({state_in_s1[263], state_in_s0[263]}), .b ({new_AGEMA_signal_3428, n3584}), .c ({new_AGEMA_signal_3713, n3563}) ) ;
    xnor_HPC2 U3717 ( .a ({new_AGEMA_signal_3989, n3560}), .b ({new_AGEMA_signal_3713, n3563}), .c ({state_out_s1[256], state_out_s0[256]}) ) ;
    xnor_HPC2 U3718 ( .a ({new_AGEMA_signal_3609, n3561}), .b ({new_AGEMA_signal_3612, n3776}), .c ({new_AGEMA_signal_3990, n3562}) ) ;
    xnor_HPC2 U3719 ( .a ({new_AGEMA_signal_3990, n3562}), .b ({new_AGEMA_signal_3713, n3563}), .c ({state_out_s1[263], state_out_s0[263]}) ) ;
    xnor_HPC2 U3720 ( .a ({new_AGEMA_signal_3585, n3926}), .b ({new_AGEMA_signal_3707, n3921}), .c ({new_AGEMA_signal_3991, n3564}) ) ;
    xnor_HPC2 U3721 ( .a ({new_AGEMA_signal_3991, n3564}), .b ({new_AGEMA_signal_3713, n3563}), .c ({state_out_s1[302], state_out_s0[302]}) ) ;
    xor_HPC2 U3722 ( .a ({new_AGEMA_signal_3221, z0[62]}), .b ({state_in_s1[6], state_in_s0[6]}), .c ({new_AGEMA_signal_3429, n3573}) ) ;
    xnor_HPC2 U3723 ( .a ({new_AGEMA_signal_3429, n3573}), .b ({new_AGEMA_signal_3417, n3565}), .c ({new_AGEMA_signal_3714, n3872}) ) ;
    xnor_HPC2 U3724 ( .a ({new_AGEMA_signal_3407, n3567}), .b ({new_AGEMA_signal_3311, n3566}), .c ({new_AGEMA_signal_3715, n3773}) ) ;
    xnor_HPC2 U3725 ( .a ({new_AGEMA_signal_3714, n3872}), .b ({new_AGEMA_signal_3715, n3773}), .c ({new_AGEMA_signal_3992, n3570}) ) ;
    xnor_HPC2 U3726 ( .a ({new_AGEMA_signal_3339, n3569}), .b ({new_AGEMA_signal_3325, n3568}), .c ({new_AGEMA_signal_3716, n3760}) ) ;
    xnor_HPC2 U3727 ( .a ({new_AGEMA_signal_3992, n3570}), .b ({new_AGEMA_signal_3716, n3760}), .c ({state_out_s1[26], state_out_s0[26]}) ) ;
    xnor_HPC2 U3728 ( .a ({new_AGEMA_signal_3910, n3572}), .b ({new_AGEMA_signal_3973, n3571}), .c ({new_AGEMA_signal_4292, n3576}) ) ;
    xor_HPC2 U3729 ( .a ({new_AGEMA_signal_3043, z1[62]}), .b ({state_in_s1[262], state_in_s0[262]}), .c ({new_AGEMA_signal_3430, n3575}) ) ;
    xnor_HPC2 U3730 ( .a ({state_in_s1[70], state_in_s0[70]}), .b ({new_AGEMA_signal_3429, n3573}), .c ({new_AGEMA_signal_3717, n3574}) ) ;
    xnor_HPC2 U3731 ( .a ({new_AGEMA_signal_3430, n3575}), .b ({new_AGEMA_signal_3717, n3574}), .c ({new_AGEMA_signal_3993, n3677}) ) ;
    xnor_HPC2 U3732 ( .a ({new_AGEMA_signal_4292, n3576}), .b ({new_AGEMA_signal_3993, n3677}), .c ({state_out_s1[70], state_out_s0[70]}) ) ;
    xnor_HPC2 U3733 ( .a ({new_AGEMA_signal_3925, n3796}), .b ({new_AGEMA_signal_3993, n3677}), .c ({new_AGEMA_signal_4293, n3579}) ) ;
    xor_HPC2 U3734 ( .a ({new_AGEMA_signal_3004, z1[23]}), .b ({state_in_s1[303], state_in_s0[303]}), .c ({new_AGEMA_signal_3431, n3578}) ) ;
    xor_HPC2 U3735 ( .a ({new_AGEMA_signal_3241, z0[23]}), .b ({state_in_s1[47], state_in_s0[47]}), .c ({new_AGEMA_signal_3432, n3595}) ) ;
    xnor_HPC2 U3736 ( .a ({state_in_s1[111], state_in_s0[111]}), .b ({new_AGEMA_signal_3432, n3595}), .c ({new_AGEMA_signal_3718, n3577}) ) ;
    xnor_HPC2 U3737 ( .a ({new_AGEMA_signal_3431, n3578}), .b ({new_AGEMA_signal_3718, n3577}), .c ({new_AGEMA_signal_3994, n3790}) ) ;
    xnor_HPC2 U3738 ( .a ({new_AGEMA_signal_4293, n3579}), .b ({new_AGEMA_signal_3994, n3790}), .c ({state_out_s1[111], state_out_s0[111]}) ) ;
    xnor_HPC2 U3739 ( .a ({new_AGEMA_signal_3350, n3581}), .b ({new_AGEMA_signal_3326, n3580}), .c ({new_AGEMA_signal_3719, n3876}) ) ;
    xnor_HPC2 U3740 ( .a ({new_AGEMA_signal_3419, n3583}), .b ({new_AGEMA_signal_3316, n3582}), .c ({new_AGEMA_signal_3720, n3859}) ) ;
    xnor_HPC2 U3741 ( .a ({new_AGEMA_signal_3719, n3876}), .b ({new_AGEMA_signal_3720, n3859}), .c ({new_AGEMA_signal_3995, n3585}) ) ;
    xor_HPC2 U3742 ( .a ({new_AGEMA_signal_3218, z0[63]}), .b ({state_in_s1[7], state_in_s0[7]}), .c ({new_AGEMA_signal_3433, n3587}) ) ;
    xnor_HPC2 U3743 ( .a ({new_AGEMA_signal_3433, n3587}), .b ({new_AGEMA_signal_3428, n3584}), .c ({new_AGEMA_signal_3721, n3855}) ) ;
    xnor_HPC2 U3744 ( .a ({new_AGEMA_signal_3995, n3585}), .b ({new_AGEMA_signal_3721, n3855}), .c ({state_out_s1[27], state_out_s0[27]}) ) ;
    xnor_HPC2 U3745 ( .a ({new_AGEMA_signal_3916, n3586}), .b ({new_AGEMA_signal_3951, n3607}), .c ({new_AGEMA_signal_4295, n3590}) ) ;
    xor_HPC2 U3746 ( .a ({new_AGEMA_signal_3044, z1[63]}), .b ({state_in_s1[263], state_in_s0[263]}), .c ({new_AGEMA_signal_3434, n3589}) ) ;
    xnor_HPC2 U3747 ( .a ({state_in_s1[71], state_in_s0[71]}), .b ({new_AGEMA_signal_3433, n3587}), .c ({new_AGEMA_signal_3722, n3588}) ) ;
    xnor_HPC2 U3748 ( .a ({new_AGEMA_signal_3434, n3589}), .b ({new_AGEMA_signal_3722, n3588}), .c ({new_AGEMA_signal_3996, n3720}) ) ;
    xnor_HPC2 U3749 ( .a ({new_AGEMA_signal_4295, n3590}), .b ({new_AGEMA_signal_3996, n3720}), .c ({state_out_s1[71], state_out_s0[71]}) ) ;
    xnor_HPC2 U3750 ( .a ({new_AGEMA_signal_3919, n3853}), .b ({new_AGEMA_signal_3996, n3720}), .c ({new_AGEMA_signal_4296, n3594}) ) ;
    xor_HPC2 U3751 ( .a ({new_AGEMA_signal_3005, z1[24]}), .b ({state_in_s1[288], state_in_s0[288]}), .c ({new_AGEMA_signal_3435, n3593}) ) ;
    xnor_HPC2 U3752 ( .a ({state_in_s1[96], state_in_s0[96]}), .b ({new_AGEMA_signal_3411, n3591}), .c ({new_AGEMA_signal_3723, n3592}) ) ;
    xnor_HPC2 U3753 ( .a ({new_AGEMA_signal_3435, n3593}), .b ({new_AGEMA_signal_3723, n3592}), .c ({new_AGEMA_signal_3997, n3848}) ) ;
    xnor_HPC2 U3754 ( .a ({new_AGEMA_signal_4296, n3594}), .b ({new_AGEMA_signal_3997, n3848}), .c ({state_out_s1[96], state_out_s0[96]}) ) ;
    xnor_HPC2 U3755 ( .a ({state_in_s1[239], state_in_s0[239]}), .b ({new_AGEMA_signal_3126, z4[23]}), .c ({new_AGEMA_signal_3436, n3601}) ) ;
    xnor_HPC2 U3756 ( .a ({new_AGEMA_signal_3432, n3595}), .b ({new_AGEMA_signal_3436, n3601}), .c ({new_AGEMA_signal_3724, n3894}) ) ;
    xnor_HPC2 U3757 ( .a ({new_AGEMA_signal_3337, n3597}), .b ({new_AGEMA_signal_3367, n3596}), .c ({new_AGEMA_signal_3725, n3890}) ) ;
    xnor_HPC2 U3758 ( .a ({new_AGEMA_signal_3724, n3894}), .b ({new_AGEMA_signal_3725, n3890}), .c ({new_AGEMA_signal_3998, n3600}) ) ;
    xnor_HPC2 U3759 ( .a ({new_AGEMA_signal_3405, n3599}), .b ({new_AGEMA_signal_3329, n3598}), .c ({new_AGEMA_signal_3726, n3737}) ) ;
    xnor_HPC2 U3760 ( .a ({new_AGEMA_signal_3998, n3600}), .b ({new_AGEMA_signal_3726, n3737}), .c ({state_out_s1[3], state_out_s0[3]}) ) ;
    xnor_HPC2 U3761 ( .a ({new_AGEMA_signal_3601, n3625}), .b ({new_AGEMA_signal_3603, n3687}), .c ({new_AGEMA_signal_3999, n3602}) ) ;
    xnor_HPC2 U3762 ( .a ({state_in_s1[303], state_in_s0[303]}), .b ({new_AGEMA_signal_3436, n3601}), .c ({new_AGEMA_signal_3727, n3690}) ) ;
    xnor_HPC2 U3763 ( .a ({new_AGEMA_signal_3999, n3602}), .b ({new_AGEMA_signal_3727, n3690}), .c ({state_out_s1[278], state_out_s0[278]}) ) ;
    xnor_HPC2 U3764 ( .a ({new_AGEMA_signal_3389, n3604}), .b ({new_AGEMA_signal_3321, n3603}), .c ({new_AGEMA_signal_3728, n3893}) ) ;
    xnor_HPC2 U3765 ( .a ({new_AGEMA_signal_3666, n3887}), .b ({new_AGEMA_signal_3728, n3893}), .c ({new_AGEMA_signal_4000, n3606}) ) ;
    xor_HPC2 U3766 ( .a ({new_AGEMA_signal_3219, z0[41]}), .b ({state_in_s1[17], state_in_s0[17]}), .c ({new_AGEMA_signal_3437, n3609}) ) ;
    xnor_HPC2 U3767 ( .a ({new_AGEMA_signal_3437, n3609}), .b ({new_AGEMA_signal_3324, n3605}), .c ({new_AGEMA_signal_3729, n3740}) ) ;
    xnor_HPC2 U3768 ( .a ({new_AGEMA_signal_4000, n3606}), .b ({new_AGEMA_signal_3729, n3740}), .c ({state_out_s1[53], state_out_s0[53]}) ) ;
    xnor_HPC2 U3769 ( .a ({new_AGEMA_signal_3922, n3608}), .b ({new_AGEMA_signal_3951, n3607}), .c ({new_AGEMA_signal_4300, n3612}) ) ;
    xor_HPC2 U3770 ( .a ({new_AGEMA_signal_3022, z1[41]}), .b ({new_AGEMA_signal_3437, n3609}), .c ({new_AGEMA_signal_3730, n3611}) ) ;
    xnor_HPC2 U3772 ( .a ({new_AGEMA_signal_3730, n3611}), .b ({new_AGEMA_signal_2685, n3610}), .c ({new_AGEMA_signal_4001, n3719}) ) ;
    xnor_HPC2 U3773 ( .a ({new_AGEMA_signal_4300, n3612}), .b ({new_AGEMA_signal_4001, n3719}), .c ({state_out_s1[81], state_out_s0[81]}) ) ;
    xnor_HPC2 U3774 ( .a ({new_AGEMA_signal_3334, n3614}), .b ({new_AGEMA_signal_3323, n3613}), .c ({new_AGEMA_signal_3731, n3915}) ) ;
    xnor_HPC2 U3775 ( .a ({new_AGEMA_signal_3726, n3737}), .b ({new_AGEMA_signal_3731, n3915}), .c ({new_AGEMA_signal_4002, n3616}) ) ;
    xor_HPC2 U3776 ( .a ({new_AGEMA_signal_3217, z0[42]}), .b ({state_in_s1[18], state_in_s0[18]}), .c ({new_AGEMA_signal_3438, n3618}) ) ;
    xnor_HPC2 U3777 ( .a ({new_AGEMA_signal_3438, n3618}), .b ({new_AGEMA_signal_3299, n3615}), .c ({new_AGEMA_signal_3732, n3828}) ) ;
    xnor_HPC2 U3778 ( .a ({new_AGEMA_signal_4002, n3616}), .b ({new_AGEMA_signal_3732, n3828}), .c ({state_out_s1[54], state_out_s0[54]}) ) ;
    xnor_HPC2 U3779 ( .a ({new_AGEMA_signal_3926, n3617}), .b ({new_AGEMA_signal_3981, n3644}), .c ({new_AGEMA_signal_4302, n3621}) ) ;
    xor_HPC2 U3780 ( .a ({new_AGEMA_signal_3023, z1[42]}), .b ({state_in_s1[274], state_in_s0[274]}), .c ({new_AGEMA_signal_3439, n3620}) ) ;
    xnor_HPC2 U3781 ( .a ({state_in_s1[82], state_in_s0[82]}), .b ({new_AGEMA_signal_3438, n3618}), .c ({new_AGEMA_signal_3733, n3619}) ) ;
    xnor_HPC2 U3782 ( .a ({new_AGEMA_signal_3439, n3620}), .b ({new_AGEMA_signal_3733, n3619}), .c ({new_AGEMA_signal_4003, n3816}) ) ;
    xnor_HPC2 U3783 ( .a ({new_AGEMA_signal_4302, n3621}), .b ({new_AGEMA_signal_4003, n3816}), .c ({state_out_s1[82], state_out_s0[82]}) ) ;
    xnor_HPC2 U3784 ( .a ({new_AGEMA_signal_3678, n3704}), .b ({new_AGEMA_signal_3703, n3802}), .c ({new_AGEMA_signal_4004, n3623}) ) ;
    xnor_HPC2 U3785 ( .a ({state_in_s1[230], state_in_s0[230]}), .b ({new_AGEMA_signal_3134, z4[30]}), .c ({new_AGEMA_signal_3440, n3626}) ) ;
    xnor_HPC2 U3786 ( .a ({new_AGEMA_signal_3371, n3622}), .b ({new_AGEMA_signal_3440, n3626}), .c ({new_AGEMA_signal_3734, n3711}) ) ;
    xnor_HPC2 U3787 ( .a ({new_AGEMA_signal_4004, n3623}), .b ({new_AGEMA_signal_3734, n3711}), .c ({state_out_s1[51], state_out_s0[51]}) ) ;
    xnor_HPC2 U3788 ( .a ({new_AGEMA_signal_3601, n3625}), .b ({new_AGEMA_signal_3661, n3624}), .c ({new_AGEMA_signal_4005, n3627}) ) ;
    xnor_HPC2 U3789 ( .a ({state_in_s1[294], state_in_s0[294]}), .b ({new_AGEMA_signal_3440, n3626}), .c ({new_AGEMA_signal_3735, n3632}) ) ;
    xnor_HPC2 U3790 ( .a ({new_AGEMA_signal_4005, n3627}), .b ({new_AGEMA_signal_3735, n3632}), .c ({state_out_s1[269], state_out_s0[269]}) ) ;
    xnor_HPC2 U3791 ( .a ({new_AGEMA_signal_3618, n3629}), .b ({new_AGEMA_signal_3655, n3628}), .c ({new_AGEMA_signal_4006, n3630}) ) ;
    xnor_HPC2 U3792 ( .a ({new_AGEMA_signal_4006, n3630}), .b ({new_AGEMA_signal_3735, n3632}), .c ({state_out_s1[294], state_out_s0[294]}) ) ;
    xnor_HPC2 U3793 ( .a ({new_AGEMA_signal_3631, n3631}), .b ({new_AGEMA_signal_3727, n3690}), .c ({new_AGEMA_signal_4007, n3633}) ) ;
    xnor_HPC2 U3794 ( .a ({new_AGEMA_signal_4007, n3633}), .b ({new_AGEMA_signal_3735, n3632}), .c ({state_out_s1[303], state_out_s0[303]}) ) ;
    xnor_HPC2 U3795 ( .a ({new_AGEMA_signal_3662, n3846}), .b ({new_AGEMA_signal_3672, n3787}), .c ({new_AGEMA_signal_4008, n3635}) ) ;
    xor_HPC2 U3796 ( .a ({new_AGEMA_signal_3584, z0[0]}), .b ({state_in_s1[56], state_in_s0[56]}), .c ({new_AGEMA_signal_3736, n3639}) ) ;
    xnor_HPC2 U3797 ( .a ({new_AGEMA_signal_3736, n3639}), .b ({new_AGEMA_signal_3345, n3634}), .c ({new_AGEMA_signal_4009, n3782}) ) ;
    xnor_HPC2 U3798 ( .a ({new_AGEMA_signal_4008, n3635}), .b ({new_AGEMA_signal_4009, n3782}), .c ({state_out_s1[28], state_out_s0[28]}) ) ;
    xnor_HPC2 U3799 ( .a ({new_AGEMA_signal_3645, n3637}), .b ({new_AGEMA_signal_3687, n3636}), .c ({new_AGEMA_signal_4010, n3638}) ) ;
    xnor_HPC2 U3800 ( .a ({new_AGEMA_signal_4010, n3638}), .b ({new_AGEMA_signal_4009, n3782}), .c ({state_out_s1[56], state_out_s0[56]}) ) ;
    xnor_HPC2 U3801 ( .a ({new_AGEMA_signal_3934, n3810}), .b ({new_AGEMA_signal_3986, n3702}), .c ({new_AGEMA_signal_4309, n3642}) ) ;
    xor_HPC2 U3802 ( .a ({new_AGEMA_signal_3517, z1[0]}), .b ({state_in_s1[312], state_in_s0[312]}), .c ({new_AGEMA_signal_3737, n3641}) ) ;
    xnor_HPC2 U3803 ( .a ({state_in_s1[120], state_in_s0[120]}), .b ({new_AGEMA_signal_3736, n3639}), .c ({new_AGEMA_signal_4011, n3640}) ) ;
    xnor_HPC2 U3804 ( .a ({new_AGEMA_signal_3737, n3641}), .b ({new_AGEMA_signal_4011, n3640}), .c ({new_AGEMA_signal_4310, n3815}) ) ;
    xnor_HPC2 U3805 ( .a ({new_AGEMA_signal_4309, n3642}), .b ({new_AGEMA_signal_4310, n3815}), .c ({state_out_s1[97], state_out_s0[97]}) ) ;
    xnor_HPC2 U3806 ( .a ({new_AGEMA_signal_3981, n3644}), .b ({new_AGEMA_signal_3985, n3643}), .c ({new_AGEMA_signal_4311, n3645}) ) ;
    xnor_HPC2 U3807 ( .a ({new_AGEMA_signal_4311, n3645}), .b ({new_AGEMA_signal_4310, n3815}), .c ({state_out_s1[120], state_out_s0[120]}) ) ;
    xnor_HPC2 U3808 ( .a ({new_AGEMA_signal_3693, n3823}), .b ({new_AGEMA_signal_3716, n3760}), .c ({new_AGEMA_signal_4012, n3647}) ) ;
    xor_HPC2 U3809 ( .a ({new_AGEMA_signal_3216, z0[43]}), .b ({state_in_s1[19], state_in_s0[19]}), .c ({new_AGEMA_signal_3441, n3649}) ) ;
    xnor_HPC2 U3810 ( .a ({new_AGEMA_signal_3441, n3649}), .b ({new_AGEMA_signal_3302, n3646}), .c ({new_AGEMA_signal_3738, n3917}) ) ;
    xnor_HPC2 U3811 ( .a ({new_AGEMA_signal_4012, n3647}), .b ({new_AGEMA_signal_3738, n3917}), .c ({state_out_s1[55], state_out_s0[55]}) ) ;
    xnor_HPC2 U3812 ( .a ({new_AGEMA_signal_3920, n3648}), .b ({new_AGEMA_signal_3988, n3678}), .c ({new_AGEMA_signal_4313, n3652}) ) ;
    xor_HPC2 U3813 ( .a ({new_AGEMA_signal_3024, z1[43]}), .b ({state_in_s1[275], state_in_s0[275]}), .c ({new_AGEMA_signal_3442, n3651}) ) ;
    xnor_HPC2 U3814 ( .a ({state_in_s1[83], state_in_s0[83]}), .b ({new_AGEMA_signal_3441, n3649}), .c ({new_AGEMA_signal_3739, n3650}) ) ;
    xnor_HPC2 U3815 ( .a ({new_AGEMA_signal_3442, n3651}), .b ({new_AGEMA_signal_3739, n3650}), .c ({new_AGEMA_signal_4013, n3904}) ) ;
    xnor_HPC2 U3816 ( .a ({new_AGEMA_signal_4313, n3652}), .b ({new_AGEMA_signal_4013, n3904}), .c ({state_out_s1[83], state_out_s0[83]}) ) ;
    xnor_HPC2 U3817 ( .a ({new_AGEMA_signal_3668, n3803}), .b ({new_AGEMA_signal_3734, n3711}), .c ({new_AGEMA_signal_4014, n3654}) ) ;
    xnor_HPC2 U3818 ( .a ({state_in_s1[201], state_in_s0[201]}), .b ({new_AGEMA_signal_3154, z4[49]}), .c ({new_AGEMA_signal_3443, n3658}) ) ;
    xnor_HPC2 U3819 ( .a ({new_AGEMA_signal_3398, n3653}), .b ({new_AGEMA_signal_3443, n3658}), .c ({new_AGEMA_signal_3740, n3886}) ) ;
    xnor_HPC2 U3820 ( .a ({new_AGEMA_signal_4014, n3654}), .b ({new_AGEMA_signal_3740, n3886}), .c ({state_out_s1[38], state_out_s0[38]}) ) ;
    xnor_HPC2 U3821 ( .a ({new_AGEMA_signal_3696, n3712}), .b ({new_AGEMA_signal_3710, n3891}), .c ({new_AGEMA_signal_4015, n3655}) ) ;
    xnor_HPC2 U3822 ( .a ({new_AGEMA_signal_4015, n3655}), .b ({new_AGEMA_signal_3740, n3886}), .c ({state_out_s1[45], state_out_s0[45]}) ) ;
    xnor_HPC2 U3823 ( .a ({new_AGEMA_signal_3587, n3657}), .b ({new_AGEMA_signal_3654, n3656}), .c ({new_AGEMA_signal_4016, n3659}) ) ;
    xnor_HPC2 U3824 ( .a ({state_in_s1[265], state_in_s0[265]}), .b ({new_AGEMA_signal_3443, n3658}), .c ({new_AGEMA_signal_3741, n3665}) ) ;
    xnor_HPC2 U3825 ( .a ({new_AGEMA_signal_4016, n3659}), .b ({new_AGEMA_signal_3741, n3665}), .c ({state_out_s1[265], state_out_s0[265]}) ) ;
    xnor_HPC2 U3826 ( .a ({new_AGEMA_signal_3589, n3661}), .b ({new_AGEMA_signal_3600, n3660}), .c ({new_AGEMA_signal_4017, n3662}) ) ;
    xnor_HPC2 U3827 ( .a ({new_AGEMA_signal_4017, n3662}), .b ({new_AGEMA_signal_3741, n3665}), .c ({state_out_s1[274], state_out_s0[274]}) ) ;
    xnor_HPC2 U3828 ( .a ({new_AGEMA_signal_3586, n3664}), .b ({new_AGEMA_signal_3588, n3663}), .c ({new_AGEMA_signal_4018, n3666}) ) ;
    xnor_HPC2 U3829 ( .a ({new_AGEMA_signal_4018, n3666}), .b ({new_AGEMA_signal_3741, n3665}), .c ({state_out_s1[304], state_out_s0[304]}) ) ;
    xnor_HPC2 U3830 ( .a ({new_AGEMA_signal_3680, n3667}), .b ({new_AGEMA_signal_3688, n3863}), .c ({new_AGEMA_signal_4019, n3669}) ) ;
    xor_HPC2 U3831 ( .a ({new_AGEMA_signal_3890, z0[1]}), .b ({state_in_s1[57], state_in_s0[57]}), .c ({new_AGEMA_signal_4020, n3673}) ) ;
    xnor_HPC2 U3832 ( .a ({new_AGEMA_signal_4020, n3673}), .b ({new_AGEMA_signal_3300, n3668}), .c ({new_AGEMA_signal_4319, n3842}) ) ;
    xnor_HPC2 U3833 ( .a ({new_AGEMA_signal_4019, n3669}), .b ({new_AGEMA_signal_4319, n3842}), .c ({state_out_s1[29], state_out_s0[29]}) ) ;
    xnor_HPC2 U3834 ( .a ({new_AGEMA_signal_3679, n3671}), .b ({new_AGEMA_signal_3706, n3670}), .c ({new_AGEMA_signal_4021, n3672}) ) ;
    xnor_HPC2 U3835 ( .a ({new_AGEMA_signal_4021, n3672}), .b ({new_AGEMA_signal_4319, n3842}), .c ({state_out_s1[57], state_out_s0[57]}) ) ;
    xnor_HPC2 U3836 ( .a ({new_AGEMA_signal_3942, n3898}), .b ({new_AGEMA_signal_3994, n3790}), .c ({new_AGEMA_signal_4320, n3676}) ) ;
    xor_HPC2 U3837 ( .a ({new_AGEMA_signal_3887, z1[1]}), .b ({state_in_s1[313], state_in_s0[313]}), .c ({new_AGEMA_signal_4022, n3675}) ) ;
    xnor_HPC2 U3838 ( .a ({state_in_s1[121], state_in_s0[121]}), .b ({new_AGEMA_signal_4020, n3673}), .c ({new_AGEMA_signal_4321, n3674}) ) ;
    xnor_HPC2 U3839 ( .a ({new_AGEMA_signal_4022, n3675}), .b ({new_AGEMA_signal_4321, n3674}), .c ({new_AGEMA_signal_4496, n3903}) ) ;
    xnor_HPC2 U3840 ( .a ({new_AGEMA_signal_4320, n3676}), .b ({new_AGEMA_signal_4496, n3903}), .c ({state_out_s1[98], state_out_s0[98]}) ) ;
    xnor_HPC2 U3841 ( .a ({new_AGEMA_signal_3988, n3678}), .b ({new_AGEMA_signal_3993, n3677}), .c ({new_AGEMA_signal_4322, n3679}) ) ;
    xnor_HPC2 U3842 ( .a ({new_AGEMA_signal_4322, n3679}), .b ({new_AGEMA_signal_4496, n3903}), .c ({state_out_s1[121], state_out_s0[121]}) ) ;
    xnor_HPC2 U3843 ( .a ({new_AGEMA_signal_3425, n3681}), .b ({new_AGEMA_signal_3403, n3680}), .c ({new_AGEMA_signal_3742, n3914}) ) ;
    xnor_HPC2 U3844 ( .a ({state_in_s1[232], state_in_s0[232]}), .b ({new_AGEMA_signal_3118, z4[16]}), .c ({new_AGEMA_signal_3444, n3688}) ) ;
    xnor_HPC2 U3845 ( .a ({new_AGEMA_signal_3357, n3682}), .b ({new_AGEMA_signal_3444, n3688}), .c ({new_AGEMA_signal_3743, n3911}) ) ;
    xnor_HPC2 U3846 ( .a ({new_AGEMA_signal_3742, n3914}), .b ({new_AGEMA_signal_3743, n3911}), .c ({new_AGEMA_signal_4023, n3685}) ) ;
    xnor_HPC2 U3847 ( .a ({new_AGEMA_signal_3372, n3684}), .b ({new_AGEMA_signal_3365, n3683}), .c ({new_AGEMA_signal_3744, n3759}) ) ;
    xnor_HPC2 U3848 ( .a ({new_AGEMA_signal_4023, n3685}), .b ({new_AGEMA_signal_3744, n3759}), .c ({state_out_s1[5], state_out_s0[5]}) ) ;
    xnor_HPC2 U3849 ( .a ({new_AGEMA_signal_3603, n3687}), .b ({new_AGEMA_signal_3610, n3686}), .c ({new_AGEMA_signal_4024, n3689}) ) ;
    xnor_HPC2 U3850 ( .a ({state_in_s1[296], state_in_s0[296]}), .b ({new_AGEMA_signal_3444, n3688}), .c ({new_AGEMA_signal_3745, n3732}) ) ;
    xnor_HPC2 U3851 ( .a ({new_AGEMA_signal_4024, n3689}), .b ({new_AGEMA_signal_3745, n3732}), .c ({state_out_s1[287], state_out_s0[287]}) ) ;
    xnor_HPC2 U3852 ( .a ({new_AGEMA_signal_3630, n3726}), .b ({new_AGEMA_signal_3727, n3690}), .c ({new_AGEMA_signal_4025, n3691}) ) ;
    xnor_HPC2 U3853 ( .a ({new_AGEMA_signal_4025, n3691}), .b ({new_AGEMA_signal_3745, n3732}), .c ({state_out_s1[296], state_out_s0[296]}) ) ;
    xnor_HPC2 U3854 ( .a ({new_AGEMA_signal_3673, n3774}), .b ({new_AGEMA_signal_3721, n3855}), .c ({new_AGEMA_signal_4026, n3693}) ) ;
    xor_HPC2 U3855 ( .a ({new_AGEMA_signal_3215, z0[44]}), .b ({state_in_s1[20], state_in_s0[20]}), .c ({new_AGEMA_signal_3445, n3698}) ) ;
    xnor_HPC2 U3856 ( .a ({new_AGEMA_signal_3445, n3698}), .b ({new_AGEMA_signal_3305, n3692}), .c ({new_AGEMA_signal_3746, n3695}) ) ;
    xnor_HPC2 U3857 ( .a ({new_AGEMA_signal_4026, n3693}), .b ({new_AGEMA_signal_3746, n3695}), .c ({state_out_s1[20], state_out_s0[20]}) ) ;
    xnor_HPC2 U3858 ( .a ({new_AGEMA_signal_3715, n3773}), .b ({new_AGEMA_signal_3744, n3759}), .c ({new_AGEMA_signal_4027, n3694}) ) ;
    xnor_HPC2 U3859 ( .a ({new_AGEMA_signal_4027, n3694}), .b ({new_AGEMA_signal_3746, n3695}), .c ({state_out_s1[33], state_out_s0[33]}) ) ;
    xnor_HPC2 U3860 ( .a ({new_AGEMA_signal_3719, n3876}), .b ({new_AGEMA_signal_3743, n3911}), .c ({new_AGEMA_signal_4028, n3696}) ) ;
    xnor_HPC2 U3861 ( .a ({new_AGEMA_signal_4028, n3696}), .b ({new_AGEMA_signal_3746, n3695}), .c ({state_out_s1[40], state_out_s0[40]}) ) ;
    xnor_HPC2 U3862 ( .a ({new_AGEMA_signal_3921, n3697}), .b ({new_AGEMA_signal_4001, n3719}), .c ({new_AGEMA_signal_4329, n3701}) ) ;
    xor_HPC2 U3863 ( .a ({new_AGEMA_signal_3025, z1[44]}), .b ({new_AGEMA_signal_3445, n3698}), .c ({new_AGEMA_signal_3747, n3700}) ) ;
    xnor_HPC2 U3865 ( .a ({new_AGEMA_signal_3747, n3700}), .b ({new_AGEMA_signal_2687, n3699}), .c ({new_AGEMA_signal_4029, n3754}) ) ;
    xnor_HPC2 U3866 ( .a ({new_AGEMA_signal_4329, n3701}), .b ({new_AGEMA_signal_4029, n3754}), .c ({state_out_s1[84], state_out_s0[84]}) ) ;
    xnor_HPC2 U3867 ( .a ({new_AGEMA_signal_3935, n3750}), .b ({new_AGEMA_signal_3986, n3702}), .c ({new_AGEMA_signal_4330, n3703}) ) ;
    xnor_HPC2 U3868 ( .a ({new_AGEMA_signal_4330, n3703}), .b ({new_AGEMA_signal_4029, n3754}), .c ({state_out_s1[87], state_out_s0[87]}) ) ;
    xnor_HPC2 U3869 ( .a ({new_AGEMA_signal_3644, n3705}), .b ({new_AGEMA_signal_3678, n3704}), .c ({new_AGEMA_signal_4030, n3707}) ) ;
    xor_HPC2 U3870 ( .a ({new_AGEMA_signal_4203, z0[2]}), .b ({state_in_s1[58], state_in_s0[58]}), .c ({new_AGEMA_signal_4331, n3715}) ) ;
    xnor_HPC2 U3871 ( .a ({new_AGEMA_signal_4331, n3715}), .b ({new_AGEMA_signal_3303, n3706}), .c ({new_AGEMA_signal_4499, n3713}) ) ;
    xnor_HPC2 U3872 ( .a ({new_AGEMA_signal_4030, n3707}), .b ({new_AGEMA_signal_4499, n3713}), .c ({state_out_s1[23], state_out_s0[23]}) ) ;
    xnor_HPC2 U3873 ( .a ({new_AGEMA_signal_3643, n3709}), .b ({new_AGEMA_signal_3697, n3708}), .c ({new_AGEMA_signal_4031, n3710}) ) ;
    xnor_HPC2 U3874 ( .a ({new_AGEMA_signal_4031, n3710}), .b ({new_AGEMA_signal_4499, n3713}), .c ({state_out_s1[30], state_out_s0[30]}) ) ;
    xnor_HPC2 U3875 ( .a ({new_AGEMA_signal_3696, n3712}), .b ({new_AGEMA_signal_3734, n3711}), .c ({new_AGEMA_signal_4032, n3714}) ) ;
    xnor_HPC2 U3876 ( .a ({new_AGEMA_signal_4032, n3714}), .b ({new_AGEMA_signal_4499, n3713}), .c ({state_out_s1[58], state_out_s0[58]}) ) ;
    xnor_HPC2 U3877 ( .a ({new_AGEMA_signal_3956, n3744}), .b ({new_AGEMA_signal_3997, n3848}), .c ({new_AGEMA_signal_4332, n3718}) ) ;
    xor_HPC2 U3878 ( .a ({new_AGEMA_signal_4200, z1[2]}), .b ({state_in_s1[314], state_in_s0[314]}), .c ({new_AGEMA_signal_4333, n3717}) ) ;
    xnor_HPC2 U3879 ( .a ({state_in_s1[122], state_in_s0[122]}), .b ({new_AGEMA_signal_4331, n3715}), .c ({new_AGEMA_signal_4500, n3716}) ) ;
    xnor_HPC2 U3880 ( .a ({new_AGEMA_signal_4333, n3717}), .b ({new_AGEMA_signal_4500, n3716}), .c ({new_AGEMA_signal_4586, n3753}) ) ;
    xnor_HPC2 U3881 ( .a ({new_AGEMA_signal_4332, n3718}), .b ({new_AGEMA_signal_4586, n3753}), .c ({state_out_s1[99], state_out_s0[99]}) ) ;
    xnor_HPC2 U3882 ( .a ({new_AGEMA_signal_3996, n3720}), .b ({new_AGEMA_signal_4001, n3719}), .c ({new_AGEMA_signal_4334, n3721}) ) ;
    xnor_HPC2 U3883 ( .a ({new_AGEMA_signal_4334, n3721}), .b ({new_AGEMA_signal_4586, n3753}), .c ({state_out_s1[122], state_out_s0[122]}) ) ;
    xnor_HPC2 U3884 ( .a ({new_AGEMA_signal_3711, n3805}), .b ({new_AGEMA_signal_3725, n3890}), .c ({new_AGEMA_signal_4033, n3723}) ) ;
    xnor_HPC2 U3885 ( .a ({state_in_s1[202], state_in_s0[202]}), .b ({new_AGEMA_signal_3156, z4[50]}), .c ({new_AGEMA_signal_3446, n3727}) ) ;
    xnor_HPC2 U3886 ( .a ({new_AGEMA_signal_3374, n3722}), .b ({new_AGEMA_signal_3446, n3727}), .c ({new_AGEMA_signal_3748, n3736}) ) ;
    xnor_HPC2 U3887 ( .a ({new_AGEMA_signal_4033, n3723}), .b ({new_AGEMA_signal_3748, n3736}), .c ({state_out_s1[39], state_out_s0[39]}) ) ;
    xnor_HPC2 U3888 ( .a ({new_AGEMA_signal_3667, n3806}), .b ({new_AGEMA_signal_3729, n3740}), .c ({new_AGEMA_signal_4034, n3724}) ) ;
    xnor_HPC2 U3889 ( .a ({new_AGEMA_signal_4034, n3724}), .b ({new_AGEMA_signal_3748, n3736}), .c ({state_out_s1[46], state_out_s0[46]}) ) ;
    xnor_HPC2 U3890 ( .a ({new_AGEMA_signal_3630, n3726}), .b ({new_AGEMA_signal_3674, n3725}), .c ({new_AGEMA_signal_4035, n3728}) ) ;
    xnor_HPC2 U3891 ( .a ({state_in_s1[266], state_in_s0[266]}), .b ({new_AGEMA_signal_3446, n3727}), .c ({new_AGEMA_signal_3749, n3734}) ) ;
    xnor_HPC2 U3892 ( .a ({new_AGEMA_signal_4035, n3728}), .b ({new_AGEMA_signal_3749, n3734}), .c ({state_out_s1[266], state_out_s0[266]}) ) ;
    xnor_HPC2 U3893 ( .a ({new_AGEMA_signal_3592, n3730}), .b ({new_AGEMA_signal_3605, n3729}), .c ({new_AGEMA_signal_4036, n3731}) ) ;
    xnor_HPC2 U3894 ( .a ({new_AGEMA_signal_4036, n3731}), .b ({new_AGEMA_signal_3749, n3734}), .c ({state_out_s1[275], state_out_s0[275]}) ) ;
    xnor_HPC2 U3895 ( .a ({new_AGEMA_signal_3591, n3733}), .b ({new_AGEMA_signal_3745, n3732}), .c ({new_AGEMA_signal_4037, n3735}) ) ;
    xnor_HPC2 U3896 ( .a ({new_AGEMA_signal_4037, n3735}), .b ({new_AGEMA_signal_3749, n3734}), .c ({state_out_s1[305], state_out_s0[305]}) ) ;
    xnor_HPC2 U3897 ( .a ({new_AGEMA_signal_3726, n3737}), .b ({new_AGEMA_signal_3748, n3736}), .c ({new_AGEMA_signal_4038, n3739}) ) ;
    xor_HPC2 U3898 ( .a ({new_AGEMA_signal_3889, z0[5]}), .b ({state_in_s1[61], state_in_s0[61]}), .c ({new_AGEMA_signal_4039, n3746}) ) ;
    xnor_HPC2 U3899 ( .a ({new_AGEMA_signal_4039, n3746}), .b ({new_AGEMA_signal_3314, n3738}), .c ({new_AGEMA_signal_4340, n3742}) ) ;
    xnor_HPC2 U3900 ( .a ({new_AGEMA_signal_4038, n3739}), .b ({new_AGEMA_signal_4340, n3742}), .c ({state_out_s1[10], state_out_s0[10]}) ) ;
    xnor_HPC2 U3901 ( .a ({new_AGEMA_signal_3692, n3826}), .b ({new_AGEMA_signal_3729, n3740}), .c ({new_AGEMA_signal_4040, n3741}) ) ;
    xnor_HPC2 U3902 ( .a ({new_AGEMA_signal_4040, n3741}), .b ({new_AGEMA_signal_4340, n3742}), .c ({state_out_s1[17], state_out_s0[17]}) ) ;
    xnor_HPC2 U3903 ( .a ({new_AGEMA_signal_3691, n3918}), .b ({new_AGEMA_signal_3731, n3915}), .c ({new_AGEMA_signal_4041, n3743}) ) ;
    xnor_HPC2 U3904 ( .a ({new_AGEMA_signal_4041, n3743}), .b ({new_AGEMA_signal_4340, n3742}), .c ({state_out_s1[61], state_out_s0[61]}) ) ;
    xnor_HPC2 U3905 ( .a ({new_AGEMA_signal_3933, n3745}), .b ({new_AGEMA_signal_3956, n3744}), .c ({new_AGEMA_signal_4341, n3749}) ) ;
    xor_HPC2 U3906 ( .a ({new_AGEMA_signal_3888, z1[5]}), .b ({state_in_s1[317], state_in_s0[317]}), .c ({new_AGEMA_signal_4042, n3748}) ) ;
    xnor_HPC2 U3907 ( .a ({state_in_s1[125], state_in_s0[125]}), .b ({new_AGEMA_signal_4039, n3746}), .c ({new_AGEMA_signal_4342, n3747}) ) ;
    xnor_HPC2 U3908 ( .a ({new_AGEMA_signal_4042, n3748}), .b ({new_AGEMA_signal_4342, n3747}), .c ({new_AGEMA_signal_4504, n3755}) ) ;
    xnor_HPC2 U3909 ( .a ({new_AGEMA_signal_4341, n3749}), .b ({new_AGEMA_signal_4504, n3755}), .c ({state_out_s1[102], state_out_s0[102]}) ) ;
    xnor_HPC2 U3910 ( .a ({new_AGEMA_signal_3932, n3751}), .b ({new_AGEMA_signal_3935, n3750}), .c ({new_AGEMA_signal_4343, n3752}) ) ;
    xnor_HPC2 U3911 ( .a ({new_AGEMA_signal_4343, n3752}), .b ({new_AGEMA_signal_4504, n3755}), .c ({state_out_s1[112], state_out_s0[112]}) ) ;
    xnor_HPC2 U3912 ( .a ({new_AGEMA_signal_4029, n3754}), .b ({new_AGEMA_signal_4586, n3753}), .c ({new_AGEMA_signal_4614, n3756}) ) ;
    xnor_HPC2 U3913 ( .a ({new_AGEMA_signal_4614, n3756}), .b ({new_AGEMA_signal_4504, n3755}), .c ({state_out_s1[125], state_out_s0[125]}) ) ;
    xnor_HPC2 U3914 ( .a ({new_AGEMA_signal_3732, n3828}), .b ({new_AGEMA_signal_3742, n3914}), .c ({new_AGEMA_signal_4043, n3758}) ) ;
    xor_HPC2 U3915 ( .a ({new_AGEMA_signal_4202, z0[6]}), .b ({state_in_s1[62], state_in_s0[62]}), .c ({new_AGEMA_signal_4344, n3763}) ) ;
    xnor_HPC2 U3916 ( .a ({new_AGEMA_signal_4344, n3763}), .b ({new_AGEMA_signal_3319, n3757}), .c ({new_AGEMA_signal_4505, n3822}) ) ;
    xnor_HPC2 U3917 ( .a ({new_AGEMA_signal_4043, n3758}), .b ({new_AGEMA_signal_4505, n3822}), .c ({state_out_s1[18], state_out_s0[18]}) ) ;
    xnor_HPC2 U3918 ( .a ({new_AGEMA_signal_3716, n3760}), .b ({new_AGEMA_signal_3744, n3759}), .c ({new_AGEMA_signal_4044, n3761}) ) ;
    xnor_HPC2 U3919 ( .a ({new_AGEMA_signal_4044, n3761}), .b ({new_AGEMA_signal_4505, n3822}), .c ({state_out_s1[62], state_out_s0[62]}) ) ;
    xnor_HPC2 U3920 ( .a ({new_AGEMA_signal_3941, n3762}), .b ({new_AGEMA_signal_3966, n3809}), .c ({new_AGEMA_signal_4345, n3766}) ) ;
    xor_HPC2 U3921 ( .a ({new_AGEMA_signal_4201, z1[6]}), .b ({state_in_s1[318], state_in_s0[318]}), .c ({new_AGEMA_signal_4346, n3765}) ) ;
    xnor_HPC2 U3922 ( .a ({state_in_s1[126], state_in_s0[126]}), .b ({new_AGEMA_signal_4344, n3763}), .c ({new_AGEMA_signal_4506, n3764}) ) ;
    xnor_HPC2 U3923 ( .a ({new_AGEMA_signal_4346, n3765}), .b ({new_AGEMA_signal_4506, n3764}), .c ({new_AGEMA_signal_4591, n3819}) ) ;
    xnor_HPC2 U3924 ( .a ({new_AGEMA_signal_4345, n3766}), .b ({new_AGEMA_signal_4591, n3819}), .c ({state_out_s1[103], state_out_s0[103]}) ) ;
    xnor_HPC2 U3925 ( .a ({new_AGEMA_signal_3940, n3767}), .b ({new_AGEMA_signal_3943, n3791}), .c ({new_AGEMA_signal_4347, n3768}) ) ;
    xnor_HPC2 U3926 ( .a ({new_AGEMA_signal_4347, n3768}), .b ({new_AGEMA_signal_4591, n3819}), .c ({state_out_s1[113], state_out_s0[113]}) ) ;
    xnor_HPC2 U3927 ( .a ({new_AGEMA_signal_3382, n3770}), .b ({new_AGEMA_signal_3375, n3769}), .c ({new_AGEMA_signal_3750, n3875}) ) ;
    xnor_HPC2 U3928 ( .a ({new_AGEMA_signal_3714, n3872}), .b ({new_AGEMA_signal_3750, n3875}), .c ({new_AGEMA_signal_4045, n3772}) ) ;
    xnor_HPC2 U3929 ( .a ({state_in_s1[233], state_in_s0[233]}), .b ({new_AGEMA_signal_3119, z4[17]}), .c ({new_AGEMA_signal_3447, n3778}) ) ;
    xnor_HPC2 U3930 ( .a ({new_AGEMA_signal_3361, n3771}), .b ({new_AGEMA_signal_3447, n3778}), .c ({new_AGEMA_signal_3751, n3786}) ) ;
    xnor_HPC2 U3931 ( .a ({new_AGEMA_signal_4045, n3772}), .b ({new_AGEMA_signal_3751, n3786}), .c ({state_out_s1[6], state_out_s0[6]}) ) ;
    xnor_HPC2 U3932 ( .a ({new_AGEMA_signal_3673, n3774}), .b ({new_AGEMA_signal_3715, n3773}), .c ({new_AGEMA_signal_4046, n3775}) ) ;
    xnor_HPC2 U3933 ( .a ({new_AGEMA_signal_4046, n3775}), .b ({new_AGEMA_signal_3751, n3786}), .c ({state_out_s1[13], state_out_s0[13]}) ) ;
    xnor_HPC2 U3934 ( .a ({new_AGEMA_signal_3608, n3777}), .b ({new_AGEMA_signal_3612, n3776}), .c ({new_AGEMA_signal_4047, n3779}) ) ;
    xnor_HPC2 U3935 ( .a ({state_in_s1[297], state_in_s0[297]}), .b ({new_AGEMA_signal_3447, n3778}), .c ({new_AGEMA_signal_3752, n3838}) ) ;
    xnor_HPC2 U3936 ( .a ({new_AGEMA_signal_4047, n3779}), .b ({new_AGEMA_signal_3752, n3838}), .c ({state_out_s1[272], state_out_s0[272]}) ) ;
    xnor_HPC2 U3937 ( .a ({new_AGEMA_signal_3639, n3780}), .b ({new_AGEMA_signal_3642, n3832}), .c ({new_AGEMA_signal_4048, n3781}) ) ;
    xnor_HPC2 U3938 ( .a ({new_AGEMA_signal_4048, n3781}), .b ({new_AGEMA_signal_3752, n3838}), .c ({state_out_s1[297], state_out_s0[297]}) ) ;
    xnor_HPC2 U3939 ( .a ({new_AGEMA_signal_3689, n3860}), .b ({new_AGEMA_signal_4009, n3782}), .c ({new_AGEMA_signal_4352, n3784}) ) ;
    xor_HPC2 U3940 ( .a ({new_AGEMA_signal_3214, z0[45]}), .b ({state_in_s1[21], state_in_s0[21]}), .c ({new_AGEMA_signal_3448, n3792}) ) ;
    xnor_HPC2 U3941 ( .a ({new_AGEMA_signal_3448, n3792}), .b ({new_AGEMA_signal_3308, n3783}), .c ({new_AGEMA_signal_3753, n3788}) ) ;
    xnor_HPC2 U3942 ( .a ({new_AGEMA_signal_4352, n3784}), .b ({new_AGEMA_signal_3753, n3788}), .c ({state_out_s1[21], state_out_s0[21]}) ) ;
    xnor_HPC2 U3943 ( .a ({new_AGEMA_signal_3720, n3859}), .b ({new_AGEMA_signal_3750, n3875}), .c ({new_AGEMA_signal_4049, n3785}) ) ;
    xnor_HPC2 U3944 ( .a ({new_AGEMA_signal_4049, n3785}), .b ({new_AGEMA_signal_3753, n3788}), .c ({state_out_s1[34], state_out_s0[34]}) ) ;
    xnor_HPC2 U3945 ( .a ({new_AGEMA_signal_3672, n3787}), .b ({new_AGEMA_signal_3751, n3786}), .c ({new_AGEMA_signal_4050, n3789}) ) ;
    xnor_HPC2 U3946 ( .a ({new_AGEMA_signal_4050, n3789}), .b ({new_AGEMA_signal_3753, n3788}), .c ({state_out_s1[41], state_out_s0[41]}) ) ;
    xnor_HPC2 U3947 ( .a ({new_AGEMA_signal_3943, n3791}), .b ({new_AGEMA_signal_3994, n3790}), .c ({new_AGEMA_signal_4355, n3795}) ) ;
    xor_HPC2 U3948 ( .a ({new_AGEMA_signal_3026, z1[45]}), .b ({new_AGEMA_signal_3448, n3792}), .c ({new_AGEMA_signal_3754, n3794}) ) ;
    xnor_HPC2 U3950 ( .a ({new_AGEMA_signal_3754, n3794}), .b ({new_AGEMA_signal_2689, n3793}), .c ({new_AGEMA_signal_4051, n3818}) ) ;
    xnor_HPC2 U3951 ( .a ({new_AGEMA_signal_4355, n3795}), .b ({new_AGEMA_signal_4051, n3818}), .c ({state_out_s1[72], state_out_s0[72]}) ) ;
    xnor_HPC2 U3952 ( .a ({new_AGEMA_signal_3925, n3796}), .b ({new_AGEMA_signal_4003, n3816}), .c ({new_AGEMA_signal_4356, n3797}) ) ;
    xnor_HPC2 U3953 ( .a ({new_AGEMA_signal_4356, n3797}), .b ({new_AGEMA_signal_4051, n3818}), .c ({state_out_s1[85], state_out_s0[85]}) ) ;
    xnor_HPC2 U3954 ( .a ({new_AGEMA_signal_3695, n3799}), .b ({new_AGEMA_signal_3704, n3798}), .c ({new_AGEMA_signal_4052, n3801}) ) ;
    xor_HPC2 U3955 ( .a ({new_AGEMA_signal_4580, z0[3]}), .b ({state_in_s1[59], state_in_s0[59]}), .c ({new_AGEMA_signal_4592, n3811}) ) ;
    xnor_HPC2 U3956 ( .a ({new_AGEMA_signal_4592, n3811}), .b ({new_AGEMA_signal_3306, n3800}), .c ({new_AGEMA_signal_4617, n3807}) ) ;
    xnor_HPC2 U3957 ( .a ({new_AGEMA_signal_4052, n3801}), .b ({new_AGEMA_signal_4617, n3807}), .c ({state_out_s1[8], state_out_s0[8]}) ) ;
    xnor_HPC2 U3958 ( .a ({new_AGEMA_signal_3668, n3803}), .b ({new_AGEMA_signal_3703, n3802}), .c ({new_AGEMA_signal_4053, n3804}) ) ;
    xnor_HPC2 U3959 ( .a ({new_AGEMA_signal_4053, n3804}), .b ({new_AGEMA_signal_4617, n3807}), .c ({state_out_s1[31], state_out_s0[31]}) ) ;
    xnor_HPC2 U3960 ( .a ({new_AGEMA_signal_3667, n3806}), .b ({new_AGEMA_signal_3711, n3805}), .c ({new_AGEMA_signal_4054, n3808}) ) ;
    xnor_HPC2 U3961 ( .a ({new_AGEMA_signal_4054, n3808}), .b ({new_AGEMA_signal_4617, n3807}), .c ({state_out_s1[59], state_out_s0[59]}) ) ;
    xnor_HPC2 U3962 ( .a ({new_AGEMA_signal_3934, n3810}), .b ({new_AGEMA_signal_3966, n3809}), .c ({new_AGEMA_signal_4357, n3814}) ) ;
    xor_HPC2 U3963 ( .a ({new_AGEMA_signal_4577, z1[3]}), .b ({state_in_s1[315], state_in_s0[315]}), .c ({new_AGEMA_signal_4593, n3813}) ) ;
    xnor_HPC2 U3964 ( .a ({state_in_s1[123], state_in_s0[123]}), .b ({new_AGEMA_signal_4592, n3811}), .c ({new_AGEMA_signal_4618, n3812}) ) ;
    xnor_HPC2 U3965 ( .a ({new_AGEMA_signal_4593, n3813}), .b ({new_AGEMA_signal_4618, n3812}), .c ({new_AGEMA_signal_4639, n3820}) ) ;
    xnor_HPC2 U3966 ( .a ({new_AGEMA_signal_4357, n3814}), .b ({new_AGEMA_signal_4639, n3820}), .c ({state_out_s1[100], state_out_s0[100]}) ) ;
    xnor_HPC2 U3967 ( .a ({new_AGEMA_signal_4003, n3816}), .b ({new_AGEMA_signal_4310, n3815}), .c ({new_AGEMA_signal_4510, n3817}) ) ;
    xnor_HPC2 U3968 ( .a ({new_AGEMA_signal_4510, n3817}), .b ({new_AGEMA_signal_4639, n3820}), .c ({state_out_s1[123], state_out_s0[123]}) ) ;
    xnor_HPC2 U3969 ( .a ({new_AGEMA_signal_4591, n3819}), .b ({new_AGEMA_signal_4051, n3818}), .c ({new_AGEMA_signal_4619, n3821}) ) ;
    xnor_HPC2 U3970 ( .a ({new_AGEMA_signal_4619, n3821}), .b ({new_AGEMA_signal_4639, n3820}), .c ({state_out_s1[126], state_out_s0[126]}) ) ;
    xnor_HPC2 U3971 ( .a ({new_AGEMA_signal_3693, n3823}), .b ({new_AGEMA_signal_4505, n3822}), .c ({new_AGEMA_signal_4594, n3825}) ) ;
    xnor_HPC2 U3972 ( .a ({state_in_s1[203], state_in_s0[203]}), .b ({new_AGEMA_signal_3157, z4[51]}), .c ({new_AGEMA_signal_3449, n3833}) ) ;
    xnor_HPC2 U3973 ( .a ({new_AGEMA_signal_3384, n3824}), .b ({new_AGEMA_signal_3449, n3833}), .c ({new_AGEMA_signal_3755, n3829}) ) ;
    xnor_HPC2 U3974 ( .a ({new_AGEMA_signal_4594, n3825}), .b ({new_AGEMA_signal_3755, n3829}), .c ({state_out_s1[11], state_out_s0[11]}) ) ;
    xnor_HPC2 U3975 ( .a ({new_AGEMA_signal_3692, n3826}), .b ({new_AGEMA_signal_3728, n3893}), .c ({new_AGEMA_signal_4055, n3827}) ) ;
    xnor_HPC2 U3976 ( .a ({new_AGEMA_signal_4055, n3827}), .b ({new_AGEMA_signal_3755, n3829}), .c ({state_out_s1[24], state_out_s0[24]}) ) ;
    xnor_HPC2 U3977 ( .a ({new_AGEMA_signal_3724, n3894}), .b ({new_AGEMA_signal_3732, n3828}), .c ({new_AGEMA_signal_4056, n3830}) ) ;
    xnor_HPC2 U3978 ( .a ({new_AGEMA_signal_4056, n3830}), .b ({new_AGEMA_signal_3755, n3829}), .c ({state_out_s1[47], state_out_s0[47]}) ) ;
    xnor_HPC2 U3979 ( .a ({new_AGEMA_signal_3642, n3832}), .b ({new_AGEMA_signal_3690, n3831}), .c ({new_AGEMA_signal_4057, n3834}) ) ;
    xnor_HPC2 U3980 ( .a ({state_in_s1[267], state_in_s0[267]}), .b ({new_AGEMA_signal_3449, n3833}), .c ({new_AGEMA_signal_3756, n3840}) ) ;
    xnor_HPC2 U3981 ( .a ({new_AGEMA_signal_4057, n3834}), .b ({new_AGEMA_signal_3756, n3840}), .c ({state_out_s1[267], state_out_s0[267]}) ) ;
    xnor_HPC2 U3982 ( .a ({new_AGEMA_signal_3595, n3836}), .b ({new_AGEMA_signal_3620, n3835}), .c ({new_AGEMA_signal_4058, n3837}) ) ;
    xnor_HPC2 U3983 ( .a ({new_AGEMA_signal_4058, n3837}), .b ({new_AGEMA_signal_3756, n3840}), .c ({state_out_s1[276], state_out_s0[276]}) ) ;
    xnor_HPC2 U3984 ( .a ({new_AGEMA_signal_3594, n3839}), .b ({new_AGEMA_signal_3752, n3838}), .c ({new_AGEMA_signal_4059, n3841}) ) ;
    xnor_HPC2 U3985 ( .a ({new_AGEMA_signal_4059, n3841}), .b ({new_AGEMA_signal_3756, n3840}), .c ({state_out_s1[306], state_out_s0[306]}) ) ;
    xnor_HPC2 U3986 ( .a ({new_AGEMA_signal_3663, n3843}), .b ({new_AGEMA_signal_4319, n3842}), .c ({new_AGEMA_signal_4511, n3845}) ) ;
    xor_HPC2 U3987 ( .a ({new_AGEMA_signal_3213, z0[46]}), .b ({state_in_s1[22], state_in_s0[22]}), .c ({new_AGEMA_signal_3450, n3849}) ) ;
    xnor_HPC2 U3988 ( .a ({new_AGEMA_signal_3450, n3849}), .b ({new_AGEMA_signal_3313, n3844}), .c ({new_AGEMA_signal_3757, n3862}) ) ;
    xnor_HPC2 U3989 ( .a ({new_AGEMA_signal_4511, n3845}), .b ({new_AGEMA_signal_3757, n3862}), .c ({state_out_s1[22], state_out_s0[22]}) ) ;
    xnor_HPC2 U3990 ( .a ({new_AGEMA_signal_3662, n3846}), .b ({new_AGEMA_signal_3671, n3856}), .c ({new_AGEMA_signal_4060, n3847}) ) ;
    xnor_HPC2 U3991 ( .a ({new_AGEMA_signal_4060, n3847}), .b ({new_AGEMA_signal_3757, n3862}), .c ({state_out_s1[35], state_out_s0[35]}) ) ;
    xnor_HPC2 U3992 ( .a ({new_AGEMA_signal_3955, n3883}), .b ({new_AGEMA_signal_3997, n3848}), .c ({new_AGEMA_signal_4364, n3852}) ) ;
    xor_HPC2 U3993 ( .a ({new_AGEMA_signal_3027, z1[46]}), .b ({state_in_s1[278], state_in_s0[278]}), .c ({new_AGEMA_signal_3451, n3851}) ) ;
    xnor_HPC2 U3994 ( .a ({state_in_s1[86], state_in_s0[86]}), .b ({new_AGEMA_signal_3450, n3849}), .c ({new_AGEMA_signal_3758, n3850}) ) ;
    xnor_HPC2 U3995 ( .a ({new_AGEMA_signal_3451, n3851}), .b ({new_AGEMA_signal_3758, n3850}), .c ({new_AGEMA_signal_4061, n3907}) ) ;
    xnor_HPC2 U3996 ( .a ({new_AGEMA_signal_4364, n3852}), .b ({new_AGEMA_signal_4061, n3907}), .c ({state_out_s1[73], state_out_s0[73]}) ) ;
    xnor_HPC2 U3997 ( .a ({new_AGEMA_signal_3919, n3853}), .b ({new_AGEMA_signal_4013, n3904}), .c ({new_AGEMA_signal_4365, n3854}) ) ;
    xnor_HPC2 U3998 ( .a ({new_AGEMA_signal_4365, n3854}), .b ({new_AGEMA_signal_4061, n3907}), .c ({state_out_s1[86], state_out_s0[86]}) ) ;
    xnor_HPC2 U3999 ( .a ({new_AGEMA_signal_3671, n3856}), .b ({new_AGEMA_signal_3721, n3855}), .c ({new_AGEMA_signal_4062, n3858}) ) ;
    xnor_HPC2 U4000 ( .a ({state_in_s1[234], state_in_s0[234]}), .b ({new_AGEMA_signal_3120, z4[18]}), .c ({new_AGEMA_signal_3452, n3868}) ) ;
    xnor_HPC2 U4001 ( .a ({new_AGEMA_signal_3353, n3857}), .b ({new_AGEMA_signal_3452, n3868}), .c ({new_AGEMA_signal_3759, n3864}) ) ;
    xnor_HPC2 U4002 ( .a ({new_AGEMA_signal_4062, n3858}), .b ({new_AGEMA_signal_3759, n3864}), .c ({state_out_s1[7], state_out_s0[7]}) ) ;
    xnor_HPC2 U4003 ( .a ({new_AGEMA_signal_3689, n3860}), .b ({new_AGEMA_signal_3720, n3859}), .c ({new_AGEMA_signal_4063, n3861}) ) ;
    xnor_HPC2 U4004 ( .a ({new_AGEMA_signal_4063, n3861}), .b ({new_AGEMA_signal_3759, n3864}), .c ({state_out_s1[14], state_out_s0[14]}) ) ;
    xnor_HPC2 U4005 ( .a ({new_AGEMA_signal_3688, n3863}), .b ({new_AGEMA_signal_3757, n3862}), .c ({new_AGEMA_signal_4064, n3865}) ) ;
    xnor_HPC2 U4006 ( .a ({new_AGEMA_signal_4064, n3865}), .b ({new_AGEMA_signal_3759, n3864}), .c ({state_out_s1[42], state_out_s0[42]}) ) ;
    xnor_HPC2 U4007 ( .a ({new_AGEMA_signal_3614, n3867}), .b ({new_AGEMA_signal_3647, n3866}), .c ({new_AGEMA_signal_4065, n3869}) ) ;
    xnor_HPC2 U4008 ( .a ({state_in_s1[298], state_in_s0[298]}), .b ({new_AGEMA_signal_3452, n3868}), .c ({new_AGEMA_signal_3760, n3928}) ) ;
    xnor_HPC2 U4009 ( .a ({new_AGEMA_signal_4065, n3869}), .b ({new_AGEMA_signal_3760, n3928}), .c ({state_out_s1[273], state_out_s0[273]}) ) ;
    xnor_HPC2 U4010 ( .a ({new_AGEMA_signal_3646, n3870}), .b ({new_AGEMA_signal_3648, n3922}), .c ({new_AGEMA_signal_4066, n3871}) ) ;
    xnor_HPC2 U4011 ( .a ({new_AGEMA_signal_4066, n3871}), .b ({new_AGEMA_signal_3760, n3928}), .c ({state_out_s1[298], state_out_s0[298]}) ) ;
    xnor_HPC2 U4012 ( .a ({new_AGEMA_signal_3714, n3872}), .b ({new_AGEMA_signal_3738, n3917}), .c ({new_AGEMA_signal_4067, n3874}) ) ;
    xor_HPC2 U4013 ( .a ({new_AGEMA_signal_4579, z0[7]}), .b ({state_in_s1[63], state_in_s0[63]}), .c ({new_AGEMA_signal_4596, n3879}) ) ;
    xnor_HPC2 U4014 ( .a ({new_AGEMA_signal_4596, n3879}), .b ({new_AGEMA_signal_3376, n3873}), .c ({new_AGEMA_signal_4621, n3910}) ) ;
    xnor_HPC2 U4015 ( .a ({new_AGEMA_signal_4067, n3874}), .b ({new_AGEMA_signal_4621, n3910}), .c ({state_out_s1[19], state_out_s0[19]}) ) ;
    xnor_HPC2 U4016 ( .a ({new_AGEMA_signal_3719, n3876}), .b ({new_AGEMA_signal_3750, n3875}), .c ({new_AGEMA_signal_4068, n3877}) ) ;
    xnor_HPC2 U4017 ( .a ({new_AGEMA_signal_4068, n3877}), .b ({new_AGEMA_signal_4621, n3910}), .c ({state_out_s1[63], state_out_s0[63]}) ) ;
    xnor_HPC2 U4018 ( .a ({new_AGEMA_signal_3949, n3878}), .b ({new_AGEMA_signal_3979, n3897}), .c ({new_AGEMA_signal_4371, n3882}) ) ;
    xor_HPC2 U4019 ( .a ({new_AGEMA_signal_4578, z1[7]}), .b ({state_in_s1[319], state_in_s0[319]}), .c ({new_AGEMA_signal_4597, n3881}) ) ;
    xnor_HPC2 U4020 ( .a ({state_in_s1[127], state_in_s0[127]}), .b ({new_AGEMA_signal_4596, n3879}), .c ({new_AGEMA_signal_4622, n3880}) ) ;
    xnor_HPC2 U4021 ( .a ({new_AGEMA_signal_4597, n3881}), .b ({new_AGEMA_signal_4622, n3880}), .c ({new_AGEMA_signal_4642, n3906}) ) ;
    xnor_HPC2 U4022 ( .a ({new_AGEMA_signal_4371, n3882}), .b ({new_AGEMA_signal_4642, n3906}), .c ({state_out_s1[88], state_out_s0[88]}) ) ;
    xnor_HPC2 U4023 ( .a ({new_AGEMA_signal_3948, n3884}), .b ({new_AGEMA_signal_3955, n3883}), .c ({new_AGEMA_signal_4372, n3885}) ) ;
    xnor_HPC2 U4024 ( .a ({new_AGEMA_signal_4372, n3885}), .b ({new_AGEMA_signal_4642, n3906}), .c ({state_out_s1[114], state_out_s0[114]}) ) ;
    xnor_HPC2 U4025 ( .a ({new_AGEMA_signal_3666, n3887}), .b ({new_AGEMA_signal_3740, n3886}), .c ({new_AGEMA_signal_4069, n3889}) ) ;
    xor_HPC2 U4026 ( .a ({new_AGEMA_signal_3583, z0[4]}), .b ({state_in_s1[60], state_in_s0[60]}), .c ({new_AGEMA_signal_3761, n3899}) ) ;
    xnor_HPC2 U4027 ( .a ({new_AGEMA_signal_3761, n3899}), .b ({new_AGEMA_signal_3309, n3888}), .c ({new_AGEMA_signal_4070, n3895}) ) ;
    xnor_HPC2 U4028 ( .a ({new_AGEMA_signal_4069, n3889}), .b ({new_AGEMA_signal_4070, n3895}), .c ({state_out_s1[9], state_out_s0[9]}) ) ;
    xnor_HPC2 U4029 ( .a ({new_AGEMA_signal_3710, n3891}), .b ({new_AGEMA_signal_3725, n3890}), .c ({new_AGEMA_signal_4071, n3892}) ) ;
    xnor_HPC2 U4030 ( .a ({new_AGEMA_signal_4071, n3892}), .b ({new_AGEMA_signal_4070, n3895}), .c ({state_out_s1[16], state_out_s0[16]}) ) ;
    xnor_HPC2 U4031 ( .a ({new_AGEMA_signal_3724, n3894}), .b ({new_AGEMA_signal_3728, n3893}), .c ({new_AGEMA_signal_4072, n3896}) ) ;
    xnor_HPC2 U4032 ( .a ({new_AGEMA_signal_4072, n3896}), .b ({new_AGEMA_signal_4070, n3895}), .c ({state_out_s1[60], state_out_s0[60]}) ) ;
    xnor_HPC2 U4033 ( .a ({new_AGEMA_signal_3942, n3898}), .b ({new_AGEMA_signal_3979, n3897}), .c ({new_AGEMA_signal_4376, n3902}) ) ;
    xor_HPC2 U4034 ( .a ({new_AGEMA_signal_3518, z1[4]}), .b ({state_in_s1[316], state_in_s0[316]}), .c ({new_AGEMA_signal_3762, n3901}) ) ;
    xnor_HPC2 U4035 ( .a ({state_in_s1[124], state_in_s0[124]}), .b ({new_AGEMA_signal_3761, n3899}), .c ({new_AGEMA_signal_4073, n3900}) ) ;
    xnor_HPC2 U4036 ( .a ({new_AGEMA_signal_3762, n3901}), .b ({new_AGEMA_signal_4073, n3900}), .c ({new_AGEMA_signal_4377, n3908}) ) ;
    xnor_HPC2 U4037 ( .a ({new_AGEMA_signal_4376, n3902}), .b ({new_AGEMA_signal_4377, n3908}), .c ({state_out_s1[101], state_out_s0[101]}) ) ;
    xnor_HPC2 U4038 ( .a ({new_AGEMA_signal_4013, n3904}), .b ({new_AGEMA_signal_4496, n3903}), .c ({new_AGEMA_signal_4598, n3905}) ) ;
    xnor_HPC2 U4039 ( .a ({new_AGEMA_signal_4598, n3905}), .b ({new_AGEMA_signal_4377, n3908}), .c ({state_out_s1[124], state_out_s0[124]}) ) ;
    xnor_HPC2 U4040 ( .a ({new_AGEMA_signal_4061, n3907}), .b ({new_AGEMA_signal_4642, n3906}), .c ({new_AGEMA_signal_4651, n3909}) ) ;
    xnor_HPC2 U4041 ( .a ({new_AGEMA_signal_4651, n3909}), .b ({new_AGEMA_signal_4377, n3908}), .c ({state_out_s1[127], state_out_s0[127]}) ) ;
    xnor_HPC2 U4042 ( .a ({new_AGEMA_signal_3743, n3911}), .b ({new_AGEMA_signal_4621, n3910}), .c ({new_AGEMA_signal_4643, n3913}) ) ;
    xnor_HPC2 U4043 ( .a ({state_in_s1[204], state_in_s0[204]}), .b ({new_AGEMA_signal_3158, z4[52]}), .c ({new_AGEMA_signal_3453, n3923}) ) ;
    xnor_HPC2 U4044 ( .a ({new_AGEMA_signal_3400, n3912}), .b ({new_AGEMA_signal_3453, n3923}), .c ({new_AGEMA_signal_3763, n3919}) ) ;
    xnor_HPC2 U4045 ( .a ({new_AGEMA_signal_4643, n3913}), .b ({new_AGEMA_signal_3763, n3919}), .c ({state_out_s1[12], state_out_s0[12]}) ) ;
    xnor_HPC2 U4046 ( .a ({new_AGEMA_signal_3731, n3915}), .b ({new_AGEMA_signal_3742, n3914}), .c ({new_AGEMA_signal_4074, n3916}) ) ;
    xnor_HPC2 U4047 ( .a ({new_AGEMA_signal_4074, n3916}), .b ({new_AGEMA_signal_3763, n3919}), .c ({state_out_s1[25], state_out_s0[25]}) ) ;
    xnor_HPC2 U4048 ( .a ({new_AGEMA_signal_3691, n3918}), .b ({new_AGEMA_signal_3738, n3917}), .c ({new_AGEMA_signal_4075, n3920}) ) ;
    xnor_HPC2 U4049 ( .a ({new_AGEMA_signal_4075, n3920}), .b ({new_AGEMA_signal_3763, n3919}), .c ({state_out_s1[32], state_out_s0[32]}) ) ;
    xnor_HPC2 U4050 ( .a ({new_AGEMA_signal_3648, n3922}), .b ({new_AGEMA_signal_3707, n3921}), .c ({new_AGEMA_signal_4076, n3924}) ) ;
    xnor_HPC2 U4051 ( .a ({state_in_s1[268], state_in_s0[268]}), .b ({new_AGEMA_signal_3453, n3923}), .c ({new_AGEMA_signal_3764, n3930}) ) ;
    xnor_HPC2 U4052 ( .a ({new_AGEMA_signal_4076, n3924}), .b ({new_AGEMA_signal_3764, n3930}), .c ({state_out_s1[268], state_out_s0[268]}) ) ;
    xnor_HPC2 U4053 ( .a ({new_AGEMA_signal_3585, n3926}), .b ({new_AGEMA_signal_3598, n3925}), .c ({new_AGEMA_signal_4077, n3927}) ) ;
    xnor_HPC2 U4054 ( .a ({new_AGEMA_signal_4077, n3927}), .b ({new_AGEMA_signal_3764, n3930}), .c ({state_out_s1[277], state_out_s0[277]}) ) ;
    xnor_HPC2 U4055 ( .a ({new_AGEMA_signal_3597, n3929}), .b ({new_AGEMA_signal_3760, n3928}), .c ({new_AGEMA_signal_4078, n3931}) ) ;
    xnor_HPC2 U4056 ( .a ({new_AGEMA_signal_4078, n3931}), .b ({new_AGEMA_signal_3764, n3930}), .c ({state_out_s1[307], state_out_s0[307]}) ) ;
    xor_HPC2 U4060 ( .a ({new_AGEMA_signal_2692, n3291}), .b ({new_AGEMA_signal_3292, z2[9]}), .c ({new_AGEMA_signal_3454, n4213}) ) ;
    xnor_HPC2 U4061 ( .a ({new_AGEMA_signal_3582, z3[9]}), .b ({state_in_s1[241], state_in_s0[241]}), .c ({new_AGEMA_signal_3765, n3932}) ) ;
    xnor_HPC2 U4062 ( .a ({new_AGEMA_signal_3454, n4213}), .b ({new_AGEMA_signal_3765, n3932}), .c ({new_AGEMA_signal_4079, n4072}) ) ;
    xor_HPC2 U4063 ( .a ({new_AGEMA_signal_2695, n3280}), .b ({new_AGEMA_signal_3282, z2[19]}), .c ({new_AGEMA_signal_3455, n4189}) ) ;
    xor_HPC2 U4064 ( .a ({new_AGEMA_signal_3529, z3[19]}), .b ({state_in_s1[235], state_in_s0[235]}), .c ({new_AGEMA_signal_3766, n3933}) ) ;
    xnor_HPC2 U4065 ( .a ({new_AGEMA_signal_3455, n4189}), .b ({new_AGEMA_signal_3766, n3933}), .c ({new_AGEMA_signal_4080, n4076}) ) ;
    xnor_HPC2 U4066 ( .a ({new_AGEMA_signal_4079, n4072}), .b ({new_AGEMA_signal_4080, n4076}), .c ({new_AGEMA_signal_4383, n3935}) ) ;
    xor_HPC2 U4067 ( .a ({new_AGEMA_signal_2698, n3273}), .b ({new_AGEMA_signal_3293, z2[26]}), .c ({new_AGEMA_signal_3456, n4174}) ) ;
    xor_HPC2 U4068 ( .a ({new_AGEMA_signal_3537, z3[26]}), .b ({state_in_s1[226], state_in_s0[226]}), .c ({new_AGEMA_signal_3767, n3934}) ) ;
    xnor_HPC2 U4069 ( .a ({new_AGEMA_signal_3456, n4174}), .b ({new_AGEMA_signal_3767, n3934}), .c ({new_AGEMA_signal_4081, n3984}) ) ;
    xnor_HPC2 U4070 ( .a ({new_AGEMA_signal_4383, n3935}), .b ({new_AGEMA_signal_4081, n3984}), .c ({state_out_s1[241], state_out_s0[241]}) ) ;
    xor_HPC2 U4074 ( .a ({new_AGEMA_signal_2701, n3279}), .b ({new_AGEMA_signal_3279, z2[20]}), .c ({new_AGEMA_signal_3457, n4186}) ) ;
    xnor_HPC2 U4075 ( .a ({new_AGEMA_signal_3531, z3[20]}), .b ({state_in_s1[236], state_in_s0[236]}), .c ({new_AGEMA_signal_3768, n3936}) ) ;
    xnor_HPC2 U4076 ( .a ({new_AGEMA_signal_3457, n4186}), .b ({new_AGEMA_signal_3768, n3936}), .c ({new_AGEMA_signal_4082, n4264}) ) ;
    xor_HPC2 U4077 ( .a ({new_AGEMA_signal_2704, n3290}), .b ({new_AGEMA_signal_3285, z2[10]}), .c ({new_AGEMA_signal_3458, n4212}) ) ;
    xor_HPC2 U4078 ( .a ({new_AGEMA_signal_3520, z3[10]}), .b ({state_in_s1[242], state_in_s0[242]}), .c ({new_AGEMA_signal_3769, n3937}) ) ;
    xnor_HPC2 U4079 ( .a ({new_AGEMA_signal_3458, n4212}), .b ({new_AGEMA_signal_3769, n3937}), .c ({new_AGEMA_signal_4083, n4269}) ) ;
    xnor_HPC2 U4080 ( .a ({new_AGEMA_signal_4082, n4264}), .b ({new_AGEMA_signal_4083, n4269}), .c ({new_AGEMA_signal_4384, n3939}) ) ;
    xor_HPC2 U4081 ( .a ({new_AGEMA_signal_2707, n3272}), .b ({new_AGEMA_signal_3291, z2[27]}), .c ({new_AGEMA_signal_3459, n4172}) ) ;
    xor_HPC2 U4082 ( .a ({new_AGEMA_signal_3538, z3[27]}), .b ({state_in_s1[227], state_in_s0[227]}), .c ({new_AGEMA_signal_3770, n3938}) ) ;
    xnor_HPC2 U4083 ( .a ({new_AGEMA_signal_3459, n4172}), .b ({new_AGEMA_signal_3770, n3938}), .c ({new_AGEMA_signal_4084, n3987}) ) ;
    xnor_HPC2 U4084 ( .a ({new_AGEMA_signal_4384, n3939}), .b ({new_AGEMA_signal_4084, n3987}), .c ({state_out_s1[242], state_out_s0[242]}) ) ;
    xor_HPC2 U4088 ( .a ({new_AGEMA_signal_2709, n3289}), .b ({new_AGEMA_signal_3283, z2[11]}), .c ({new_AGEMA_signal_3460, n4204}) ) ;
    xnor_HPC2 U4089 ( .a ({new_AGEMA_signal_3521, z3[11]}), .b ({state_in_s1[243], state_in_s0[243]}), .c ({new_AGEMA_signal_3771, n3940}) ) ;
    xnor_HPC2 U4090 ( .a ({new_AGEMA_signal_3460, n4204}), .b ({new_AGEMA_signal_3771, n3940}), .c ({new_AGEMA_signal_4085, n4258}) ) ;
    xor_HPC2 U4091 ( .a ({new_AGEMA_signal_2712, n3278}), .b ({new_AGEMA_signal_3278, z2[21]}), .c ({new_AGEMA_signal_3461, n4184}) ) ;
    xnor_HPC2 U4092 ( .a ({new_AGEMA_signal_3532, z3[21]}), .b ({state_in_s1[237], state_in_s0[237]}), .c ({new_AGEMA_signal_3772, n3941}) ) ;
    xnor_HPC2 U4093 ( .a ({new_AGEMA_signal_3461, n4184}), .b ({new_AGEMA_signal_3772, n3941}), .c ({new_AGEMA_signal_4086, n4254}) ) ;
    xor_HPC2 U4094 ( .a ({new_AGEMA_signal_2714, n3271}), .b ({new_AGEMA_signal_3290, z2[28]}), .c ({new_AGEMA_signal_3462, n4170}) ) ;
    xnor_HPC2 U4095 ( .a ({new_AGEMA_signal_3539, z3[28]}), .b ({state_in_s1[228], state_in_s0[228]}), .c ({new_AGEMA_signal_3773, n3942}) ) ;
    xnor_HPC2 U4096 ( .a ({new_AGEMA_signal_3462, n4170}), .b ({new_AGEMA_signal_3773, n3942}), .c ({new_AGEMA_signal_4087, n3989}) ) ;
    xnor_HPC2 U4097 ( .a ({new_AGEMA_signal_4086, n4254}), .b ({new_AGEMA_signal_4087, n3989}), .c ({new_AGEMA_signal_4385, n3943}) ) ;
    xnor_HPC2 U4098 ( .a ({new_AGEMA_signal_4085, n4258}), .b ({new_AGEMA_signal_4385, n3943}), .c ({state_out_s1[243], state_out_s0[243]}) ) ;
    xor_HPC2 U4102 ( .a ({new_AGEMA_signal_2717, n3288}), .b ({new_AGEMA_signal_3281, z2[12]}), .c ({new_AGEMA_signal_3463, n4192}) ) ;
    xnor_HPC2 U4103 ( .a ({new_AGEMA_signal_3522, z3[12]}), .b ({state_in_s1[244], state_in_s0[244]}), .c ({new_AGEMA_signal_3774, n3944}) ) ;
    xnor_HPC2 U4104 ( .a ({new_AGEMA_signal_3463, n4192}), .b ({new_AGEMA_signal_3774, n3944}), .c ({new_AGEMA_signal_4088, n4245}) ) ;
    xor_HPC2 U4105 ( .a ({new_AGEMA_signal_2719, n3277}), .b ({new_AGEMA_signal_3275, z2[22]}), .c ({new_AGEMA_signal_3464, n4183}) ) ;
    xnor_HPC2 U4106 ( .a ({new_AGEMA_signal_3533, z3[22]}), .b ({state_in_s1[238], state_in_s0[238]}), .c ({new_AGEMA_signal_3775, n3945}) ) ;
    xnor_HPC2 U4107 ( .a ({new_AGEMA_signal_3464, n4183}), .b ({new_AGEMA_signal_3775, n3945}), .c ({new_AGEMA_signal_4089, n4241}) ) ;
    xor_HPC2 U4108 ( .a ({new_AGEMA_signal_2721, n3270}), .b ({new_AGEMA_signal_3289, z2[29]}), .c ({new_AGEMA_signal_3465, n4169}) ) ;
    xnor_HPC2 U4109 ( .a ({new_AGEMA_signal_3540, z3[29]}), .b ({state_in_s1[229], state_in_s0[229]}), .c ({new_AGEMA_signal_3776, n3946}) ) ;
    xnor_HPC2 U4110 ( .a ({new_AGEMA_signal_3465, n4169}), .b ({new_AGEMA_signal_3776, n3946}), .c ({new_AGEMA_signal_4090, n3992}) ) ;
    xnor_HPC2 U4111 ( .a ({new_AGEMA_signal_4089, n4241}), .b ({new_AGEMA_signal_4090, n3992}), .c ({new_AGEMA_signal_4386, n3947}) ) ;
    xnor_HPC2 U4112 ( .a ({new_AGEMA_signal_4088, n4245}), .b ({new_AGEMA_signal_4386, n3947}), .c ({state_out_s1[244], state_out_s0[244]}) ) ;
    xor_HPC2 U4116 ( .a ({new_AGEMA_signal_2724, n3276}), .b ({new_AGEMA_signal_3273, z2[23]}), .c ({new_AGEMA_signal_3466, n4180}) ) ;
    xnor_HPC2 U4117 ( .a ({new_AGEMA_signal_3534, z3[23]}), .b ({state_in_s1[239], state_in_s0[239]}), .c ({new_AGEMA_signal_3777, n3948}) ) ;
    xnor_HPC2 U4118 ( .a ({new_AGEMA_signal_3466, n4180}), .b ({new_AGEMA_signal_3777, n3948}), .c ({new_AGEMA_signal_4091, n4230}) ) ;
    xor_HPC2 U4119 ( .a ({new_AGEMA_signal_2727, n3286}), .b ({new_AGEMA_signal_3280, z2[13]}), .c ({new_AGEMA_signal_3467, n4201}) ) ;
    xor_HPC2 U4120 ( .a ({new_AGEMA_signal_3523, z3[13]}), .b ({state_in_s1[245], state_in_s0[245]}), .c ({new_AGEMA_signal_3778, n3949}) ) ;
    xnor_HPC2 U4121 ( .a ({new_AGEMA_signal_3467, n4201}), .b ({new_AGEMA_signal_3778, n3949}), .c ({new_AGEMA_signal_4092, n4263}) ) ;
    xnor_HPC2 U4122 ( .a ({new_AGEMA_signal_4091, n4230}), .b ({new_AGEMA_signal_4092, n4263}), .c ({new_AGEMA_signal_4387, n3951}) ) ;
    xor_HPC2 U4123 ( .a ({new_AGEMA_signal_2730, n3269}), .b ({new_AGEMA_signal_3288, z2[30]}), .c ({new_AGEMA_signal_3468, n4166}) ) ;
    xor_HPC2 U4124 ( .a ({new_AGEMA_signal_3542, z3[30]}), .b ({state_in_s1[230], state_in_s0[230]}), .c ({new_AGEMA_signal_3779, n3950}) ) ;
    xnor_HPC2 U4125 ( .a ({new_AGEMA_signal_3468, n4166}), .b ({new_AGEMA_signal_3779, n3950}), .c ({new_AGEMA_signal_4093, n3996}) ) ;
    xnor_HPC2 U4126 ( .a ({new_AGEMA_signal_4387, n3951}), .b ({new_AGEMA_signal_4093, n3996}), .c ({state_out_s1[245], state_out_s0[245]}) ) ;
    xor_HPC2 U4130 ( .a ({new_AGEMA_signal_2733, n3285}), .b ({new_AGEMA_signal_3277, z2[14]}), .c ({new_AGEMA_signal_3469, n4199}) ) ;
    xnor_HPC2 U4131 ( .a ({new_AGEMA_signal_3524, z3[14]}), .b ({state_in_s1[246], state_in_s0[246]}), .c ({new_AGEMA_signal_3780, n3952}) ) ;
    xnor_HPC2 U4132 ( .a ({new_AGEMA_signal_3469, n4199}), .b ({new_AGEMA_signal_3780, n3952}), .c ({new_AGEMA_signal_4094, n4255}) ) ;
    xor_HPC2 U4133 ( .a ({new_AGEMA_signal_2736, n3275}), .b ({new_AGEMA_signal_3271, z2[24]}), .c ({new_AGEMA_signal_3470, n4178}) ) ;
    xnor_HPC2 U4134 ( .a ({new_AGEMA_signal_3535, z3[24]}), .b ({state_in_s1[224], state_in_s0[224]}), .c ({new_AGEMA_signal_3781, n3953}) ) ;
    xnor_HPC2 U4135 ( .a ({new_AGEMA_signal_3470, n4178}), .b ({new_AGEMA_signal_3781, n3953}), .c ({new_AGEMA_signal_4095, n4094}) ) ;
    xnor_HPC2 U4136 ( .a ({new_AGEMA_signal_4094, n4255}), .b ({new_AGEMA_signal_4095, n4094}), .c ({new_AGEMA_signal_4388, n3955}) ) ;
    xor_HPC2 U4137 ( .a ({new_AGEMA_signal_2739, n3268}), .b ({new_AGEMA_signal_3287, z2[31]}), .c ({new_AGEMA_signal_3471, n4164}) ) ;
    xnor_HPC2 U4138 ( .a ({new_AGEMA_signal_3543, z3[31]}), .b ({state_in_s1[231], state_in_s0[231]}), .c ({new_AGEMA_signal_3782, n3954}) ) ;
    xnor_HPC2 U4139 ( .a ({new_AGEMA_signal_3471, n4164}), .b ({new_AGEMA_signal_3782, n3954}), .c ({new_AGEMA_signal_4096, n3998}) ) ;
    xnor_HPC2 U4140 ( .a ({new_AGEMA_signal_4388, n3955}), .b ({new_AGEMA_signal_4096, n3998}), .c ({state_out_s1[246], state_out_s0[246]}) ) ;
    xor_HPC2 U4144 ( .a ({new_AGEMA_signal_2742, n3284}), .b ({new_AGEMA_signal_3276, z2[15]}), .c ({new_AGEMA_signal_3472, n4198}) ) ;
    xnor_HPC2 U4145 ( .a ({new_AGEMA_signal_3525, z3[15]}), .b ({state_in_s1[247], state_in_s0[247]}), .c ({new_AGEMA_signal_3783, n3956}) ) ;
    xnor_HPC2 U4146 ( .a ({new_AGEMA_signal_3472, n4198}), .b ({new_AGEMA_signal_3783, n3956}), .c ({new_AGEMA_signal_4097, n4239}) ) ;
    xor_HPC2 U4147 ( .a ({new_AGEMA_signal_2744, n3274}), .b ({new_AGEMA_signal_3286, z2[25]}), .c ({new_AGEMA_signal_3473, n4177}) ) ;
    xnor_HPC2 U4148 ( .a ({new_AGEMA_signal_3536, z3[25]}), .b ({state_in_s1[225], state_in_s0[225]}), .c ({new_AGEMA_signal_3784, n3957}) ) ;
    xnor_HPC2 U4149 ( .a ({new_AGEMA_signal_3473, n4177}), .b ({new_AGEMA_signal_3784, n3957}), .c ({new_AGEMA_signal_4098, n4044}) ) ;
    xor_HPC2 U4150 ( .a ({new_AGEMA_signal_2747, n3267}), .b ({new_AGEMA_signal_3188, z2[32]}), .c ({new_AGEMA_signal_3474, n4163}) ) ;
    xnor_HPC2 U4151 ( .a ({new_AGEMA_signal_3544, z3[32]}), .b ({state_in_s1[216], state_in_s0[216]}), .c ({new_AGEMA_signal_3785, n3958}) ) ;
    xnor_HPC2 U4152 ( .a ({new_AGEMA_signal_3474, n4163}), .b ({new_AGEMA_signal_3785, n3958}), .c ({new_AGEMA_signal_4099, n4002}) ) ;
    xnor_HPC2 U4153 ( .a ({new_AGEMA_signal_4098, n4044}), .b ({new_AGEMA_signal_4099, n4002}), .c ({new_AGEMA_signal_4389, n3959}) ) ;
    xnor_HPC2 U4154 ( .a ({new_AGEMA_signal_4097, n4239}), .b ({new_AGEMA_signal_4389, n3959}), .c ({state_out_s1[247], state_out_s0[247]}) ) ;
    xor_HPC2 U4157 ( .a ({new_AGEMA_signal_2750, n3283}), .b ({new_AGEMA_signal_3274, z2[16]}), .c ({new_AGEMA_signal_3475, n4195}) ) ;
    xnor_HPC2 U4158 ( .a ({new_AGEMA_signal_3526, z3[16]}), .b ({state_in_s1[232], state_in_s0[232]}), .c ({new_AGEMA_signal_3786, n3960}) ) ;
    xnor_HPC2 U4159 ( .a ({new_AGEMA_signal_3475, n4195}), .b ({new_AGEMA_signal_3786, n3960}), .c ({new_AGEMA_signal_4100, n4229}) ) ;
    xnor_HPC2 U4160 ( .a ({new_AGEMA_signal_4100, n4229}), .b ({new_AGEMA_signal_4081, n3984}), .c ({new_AGEMA_signal_4390, n3962}) ) ;
    xor_HPC2 U4161 ( .a ({new_AGEMA_signal_2753, n3266}), .b ({new_AGEMA_signal_3187, z2[33]}), .c ({new_AGEMA_signal_3476, n4161}) ) ;
    xor_HPC2 U4162 ( .a ({new_AGEMA_signal_3545, z3[33]}), .b ({state_in_s1[217], state_in_s0[217]}), .c ({new_AGEMA_signal_3787, n3961}) ) ;
    xnor_HPC2 U4163 ( .a ({new_AGEMA_signal_3476, n4161}), .b ({new_AGEMA_signal_3787, n3961}), .c ({new_AGEMA_signal_4101, n4006}) ) ;
    xnor_HPC2 U4164 ( .a ({new_AGEMA_signal_4390, n3962}), .b ({new_AGEMA_signal_4101, n4006}), .c ({state_out_s1[232], state_out_s0[232]}) ) ;
    xor_HPC2 U4167 ( .a ({new_AGEMA_signal_2755, n3282}), .b ({new_AGEMA_signal_3270, z2[17]}), .c ({new_AGEMA_signal_3477, n4193}) ) ;
    xnor_HPC2 U4168 ( .a ({new_AGEMA_signal_3527, z3[17]}), .b ({state_in_s1[233], state_in_s0[233]}), .c ({new_AGEMA_signal_3788, n3963}) ) ;
    xnor_HPC2 U4169 ( .a ({new_AGEMA_signal_3477, n4193}), .b ({new_AGEMA_signal_3788, n3963}), .c ({new_AGEMA_signal_4102, n4095}) ) ;
    xnor_HPC2 U4170 ( .a ({new_AGEMA_signal_4102, n4095}), .b ({new_AGEMA_signal_4084, n3987}), .c ({new_AGEMA_signal_4391, n3965}) ) ;
    xor_HPC2 U4171 ( .a ({new_AGEMA_signal_2758, n3265}), .b ({new_AGEMA_signal_3186, z2[34]}), .c ({new_AGEMA_signal_3478, n4159}) ) ;
    xor_HPC2 U4172 ( .a ({new_AGEMA_signal_3546, z3[34]}), .b ({state_in_s1[218], state_in_s0[218]}), .c ({new_AGEMA_signal_3789, n3964}) ) ;
    xnor_HPC2 U4173 ( .a ({new_AGEMA_signal_3478, n4159}), .b ({new_AGEMA_signal_3789, n3964}), .c ({new_AGEMA_signal_4103, n4007}) ) ;
    xnor_HPC2 U4174 ( .a ({new_AGEMA_signal_4391, n3965}), .b ({new_AGEMA_signal_4103, n4007}), .c ({state_out_s1[233], state_out_s0[233]}) ) ;
    xor_HPC2 U4177 ( .a ({new_AGEMA_signal_2760, n3281}), .b ({new_AGEMA_signal_3284, z2[18]}), .c ({new_AGEMA_signal_3479, n4191}) ) ;
    xnor_HPC2 U4178 ( .a ({new_AGEMA_signal_3528, z3[18]}), .b ({state_in_s1[234], state_in_s0[234]}), .c ({new_AGEMA_signal_3790, n3966}) ) ;
    xnor_HPC2 U4179 ( .a ({new_AGEMA_signal_3479, n4191}), .b ({new_AGEMA_signal_3790, n3966}), .c ({new_AGEMA_signal_4104, n4063}) ) ;
    xor_HPC2 U4180 ( .a ({new_AGEMA_signal_2763, n3264}), .b ({new_AGEMA_signal_3185, z2[35]}), .c ({new_AGEMA_signal_3480, n4157}) ) ;
    xnor_HPC2 U4181 ( .a ({new_AGEMA_signal_3547, z3[35]}), .b ({state_in_s1[219], state_in_s0[219]}), .c ({new_AGEMA_signal_3791, n3967}) ) ;
    xnor_HPC2 U4182 ( .a ({new_AGEMA_signal_3480, n4157}), .b ({new_AGEMA_signal_3791, n3967}), .c ({new_AGEMA_signal_4105, n4010}) ) ;
    xnor_HPC2 U4183 ( .a ({new_AGEMA_signal_4104, n4063}), .b ({new_AGEMA_signal_4105, n4010}), .c ({new_AGEMA_signal_4392, n3968}) ) ;
    xnor_HPC2 U4184 ( .a ({new_AGEMA_signal_4087, n3989}), .b ({new_AGEMA_signal_4392, n3968}), .c ({state_out_s1[234], state_out_s0[234]}) ) ;
    xnor_HPC2 U4186 ( .a ({new_AGEMA_signal_4090, n3992}), .b ({new_AGEMA_signal_4080, n4076}), .c ({new_AGEMA_signal_4393, n3970}) ) ;
    xor_HPC2 U4187 ( .a ({new_AGEMA_signal_2766, n3263}), .b ({new_AGEMA_signal_3183, z2[36]}), .c ({new_AGEMA_signal_3481, n4155}) ) ;
    xor_HPC2 U4188 ( .a ({new_AGEMA_signal_3548, z3[36]}), .b ({state_in_s1[220], state_in_s0[220]}), .c ({new_AGEMA_signal_3792, n3969}) ) ;
    xnor_HPC2 U4189 ( .a ({new_AGEMA_signal_3481, n4155}), .b ({new_AGEMA_signal_3792, n3969}), .c ({new_AGEMA_signal_4106, n4015}) ) ;
    xnor_HPC2 U4190 ( .a ({new_AGEMA_signal_4393, n3970}), .b ({new_AGEMA_signal_4106, n4015}), .c ({state_out_s1[235], state_out_s0[235]}) ) ;
    xnor_HPC2 U4192 ( .a ({new_AGEMA_signal_4082, n4264}), .b ({new_AGEMA_signal_4093, n3996}), .c ({new_AGEMA_signal_4394, n3972}) ) ;
    xor_HPC2 U4193 ( .a ({new_AGEMA_signal_2769, n3262}), .b ({new_AGEMA_signal_3181, z2[37]}), .c ({new_AGEMA_signal_3482, n4153}) ) ;
    xor_HPC2 U4194 ( .a ({new_AGEMA_signal_3549, z3[37]}), .b ({state_in_s1[221], state_in_s0[221]}), .c ({new_AGEMA_signal_3793, n3971}) ) ;
    xnor_HPC2 U4195 ( .a ({new_AGEMA_signal_3482, n4153}), .b ({new_AGEMA_signal_3793, n3971}), .c ({new_AGEMA_signal_4107, n4018}) ) ;
    xnor_HPC2 U4196 ( .a ({new_AGEMA_signal_4394, n3972}), .b ({new_AGEMA_signal_4107, n4018}), .c ({state_out_s1[236], state_out_s0[236]}) ) ;
    xnor_HPC2 U4198 ( .a ({new_AGEMA_signal_4086, n4254}), .b ({new_AGEMA_signal_4096, n3998}), .c ({new_AGEMA_signal_4395, n3974}) ) ;
    xor_HPC2 U4199 ( .a ({new_AGEMA_signal_2772, n3261}), .b ({new_AGEMA_signal_3179, z2[38]}), .c ({new_AGEMA_signal_3483, n4151}) ) ;
    xnor_HPC2 U4200 ( .a ({new_AGEMA_signal_3550, z3[38]}), .b ({state_in_s1[222], state_in_s0[222]}), .c ({new_AGEMA_signal_3794, n3973}) ) ;
    xnor_HPC2 U4201 ( .a ({new_AGEMA_signal_3483, n4151}), .b ({new_AGEMA_signal_3794, n3973}), .c ({new_AGEMA_signal_4108, n4019}) ) ;
    xnor_HPC2 U4202 ( .a ({new_AGEMA_signal_4395, n3974}), .b ({new_AGEMA_signal_4108, n4019}), .c ({state_out_s1[237], state_out_s0[237]}) ) ;
    xnor_HPC2 U4204 ( .a ({new_AGEMA_signal_4089, n4241}), .b ({new_AGEMA_signal_4099, n4002}), .c ({new_AGEMA_signal_4396, n3976}) ) ;
    xor_HPC2 U4205 ( .a ({new_AGEMA_signal_2775, n3260}), .b ({new_AGEMA_signal_3176, z2[39]}), .c ({new_AGEMA_signal_3484, n4149}) ) ;
    xnor_HPC2 U4206 ( .a ({new_AGEMA_signal_3551, z3[39]}), .b ({state_in_s1[223], state_in_s0[223]}), .c ({new_AGEMA_signal_3795, n3975}) ) ;
    xnor_HPC2 U4207 ( .a ({new_AGEMA_signal_3484, n4149}), .b ({new_AGEMA_signal_3795, n3975}), .c ({new_AGEMA_signal_4109, n4023}) ) ;
    xnor_HPC2 U4208 ( .a ({new_AGEMA_signal_4396, n3976}), .b ({new_AGEMA_signal_4109, n4023}), .c ({state_out_s1[238], state_out_s0[238]}) ) ;
    xnor_HPC2 U4210 ( .a ({new_AGEMA_signal_4091, n4230}), .b ({new_AGEMA_signal_4101, n4006}), .c ({new_AGEMA_signal_4397, n3978}) ) ;
    xor_HPC2 U4211 ( .a ({new_AGEMA_signal_2778, n3259}), .b ({new_AGEMA_signal_3177, z2[40]}), .c ({new_AGEMA_signal_3485, n4147}) ) ;
    xor_HPC2 U4212 ( .a ({new_AGEMA_signal_3553, z3[40]}), .b ({state_in_s1[208], state_in_s0[208]}), .c ({new_AGEMA_signal_3796, n3977}) ) ;
    xnor_HPC2 U4213 ( .a ({new_AGEMA_signal_3485, n4147}), .b ({new_AGEMA_signal_3796, n3977}), .c ({new_AGEMA_signal_4110, n4027}) ) ;
    xnor_HPC2 U4214 ( .a ({new_AGEMA_signal_4397, n3978}), .b ({new_AGEMA_signal_4110, n4027}), .c ({state_out_s1[239], state_out_s0[239]}) ) ;
    xnor_HPC2 U4216 ( .a ({new_AGEMA_signal_4095, n4094}), .b ({new_AGEMA_signal_4103, n4007}), .c ({new_AGEMA_signal_4398, n3980}) ) ;
    xor_HPC2 U4217 ( .a ({new_AGEMA_signal_2780, n3258}), .b ({new_AGEMA_signal_3184, z2[41]}), .c ({new_AGEMA_signal_3486, n4145}) ) ;
    xor_HPC2 U4218 ( .a ({new_AGEMA_signal_3554, z3[41]}), .b ({state_in_s1[209], state_in_s0[209]}), .c ({new_AGEMA_signal_3797, n3979}) ) ;
    xnor_HPC2 U4219 ( .a ({new_AGEMA_signal_3486, n4145}), .b ({new_AGEMA_signal_3797, n3979}), .c ({new_AGEMA_signal_4111, n4029}) ) ;
    xnor_HPC2 U4220 ( .a ({new_AGEMA_signal_4398, n3980}), .b ({new_AGEMA_signal_4111, n4029}), .c ({state_out_s1[224], state_out_s0[224]}) ) ;
    xnor_HPC2 U4222 ( .a ({new_AGEMA_signal_4098, n4044}), .b ({new_AGEMA_signal_4105, n4010}), .c ({new_AGEMA_signal_4399, n3982}) ) ;
    xor_HPC2 U4223 ( .a ({new_AGEMA_signal_2783, n3257}), .b ({new_AGEMA_signal_3182, z2[42]}), .c ({new_AGEMA_signal_3487, n4143}) ) ;
    xnor_HPC2 U4224 ( .a ({new_AGEMA_signal_3555, z3[42]}), .b ({state_in_s1[210], state_in_s0[210]}), .c ({new_AGEMA_signal_3798, n3981}) ) ;
    xnor_HPC2 U4225 ( .a ({new_AGEMA_signal_3487, n4143}), .b ({new_AGEMA_signal_3798, n3981}), .c ({new_AGEMA_signal_4112, n4032}) ) ;
    xnor_HPC2 U4226 ( .a ({new_AGEMA_signal_4399, n3982}), .b ({new_AGEMA_signal_4112, n4032}), .c ({state_out_s1[225], state_out_s0[225]}) ) ;
    xor_HPC2 U4228 ( .a ({new_AGEMA_signal_2786, n3256}), .b ({new_AGEMA_signal_3180, z2[43]}), .c ({new_AGEMA_signal_3488, n4141}) ) ;
    xnor_HPC2 U4229 ( .a ({new_AGEMA_signal_3556, z3[43]}), .b ({state_in_s1[211], state_in_s0[211]}), .c ({new_AGEMA_signal_3799, n3983}) ) ;
    xnor_HPC2 U4230 ( .a ({new_AGEMA_signal_3488, n4141}), .b ({new_AGEMA_signal_3799, n3983}), .c ({new_AGEMA_signal_4113, n4035}) ) ;
    xnor_HPC2 U4231 ( .a ({new_AGEMA_signal_4113, n4035}), .b ({new_AGEMA_signal_4081, n3984}), .c ({new_AGEMA_signal_4400, n3985}) ) ;
    xnor_HPC2 U4232 ( .a ({new_AGEMA_signal_4400, n3985}), .b ({new_AGEMA_signal_4106, n4015}), .c ({state_out_s1[226], state_out_s0[226]}) ) ;
    xor_HPC2 U4234 ( .a ({new_AGEMA_signal_2788, n3255}), .b ({new_AGEMA_signal_3178, z2[44]}), .c ({new_AGEMA_signal_3489, n4139}) ) ;
    xnor_HPC2 U4235 ( .a ({new_AGEMA_signal_3557, z3[44]}), .b ({state_in_s1[212], state_in_s0[212]}), .c ({new_AGEMA_signal_3800, n3986}) ) ;
    xnor_HPC2 U4236 ( .a ({new_AGEMA_signal_3489, n4139}), .b ({new_AGEMA_signal_3800, n3986}), .c ({new_AGEMA_signal_4114, n4046}) ) ;
    xnor_HPC2 U4237 ( .a ({new_AGEMA_signal_4114, n4046}), .b ({new_AGEMA_signal_4084, n3987}), .c ({new_AGEMA_signal_4401, n3988}) ) ;
    xnor_HPC2 U4238 ( .a ({new_AGEMA_signal_4401, n3988}), .b ({new_AGEMA_signal_4107, n4018}), .c ({state_out_s1[227], state_out_s0[227]}) ) ;
    xnor_HPC2 U4240 ( .a ({new_AGEMA_signal_4087, n3989}), .b ({new_AGEMA_signal_4108, n4019}), .c ({new_AGEMA_signal_4402, n3991}) ) ;
    xor_HPC2 U4241 ( .a ({new_AGEMA_signal_2790, n3254}), .b ({new_AGEMA_signal_3175, z2[45]}), .c ({new_AGEMA_signal_3490, n4137}) ) ;
    xnor_HPC2 U4242 ( .a ({new_AGEMA_signal_3558, z3[45]}), .b ({state_in_s1[213], state_in_s0[213]}), .c ({new_AGEMA_signal_3801, n3990}) ) ;
    xnor_HPC2 U4243 ( .a ({new_AGEMA_signal_3490, n4137}), .b ({new_AGEMA_signal_3801, n3990}), .c ({new_AGEMA_signal_4115, n4050}) ) ;
    xnor_HPC2 U4244 ( .a ({new_AGEMA_signal_4402, n3991}), .b ({new_AGEMA_signal_4115, n4050}), .c ({state_out_s1[228], state_out_s0[228]}) ) ;
    xnor_HPC2 U4246 ( .a ({new_AGEMA_signal_4090, n3992}), .b ({new_AGEMA_signal_4109, n4023}), .c ({new_AGEMA_signal_4403, n3994}) ) ;
    xor_HPC2 U4247 ( .a ({new_AGEMA_signal_2793, n3253}), .b ({new_AGEMA_signal_3193, z2[46]}), .c ({new_AGEMA_signal_3491, n4135}) ) ;
    xnor_HPC2 U4248 ( .a ({new_AGEMA_signal_3559, z3[46]}), .b ({state_in_s1[214], state_in_s0[214]}), .c ({new_AGEMA_signal_3802, n3993}) ) ;
    xnor_HPC2 U4249 ( .a ({new_AGEMA_signal_3491, n4135}), .b ({new_AGEMA_signal_3802, n3993}), .c ({new_AGEMA_signal_4116, n4055}) ) ;
    xnor_HPC2 U4250 ( .a ({new_AGEMA_signal_4403, n3994}), .b ({new_AGEMA_signal_4116, n4055}), .c ({state_out_s1[229], state_out_s0[229]}) ) ;
    xor_HPC2 U4252 ( .a ({new_AGEMA_signal_2795, n3252}), .b ({new_AGEMA_signal_3191, z2[47]}), .c ({new_AGEMA_signal_3492, n4133}) ) ;
    xnor_HPC2 U4253 ( .a ({new_AGEMA_signal_3560, z3[47]}), .b ({state_in_s1[215], state_in_s0[215]}), .c ({new_AGEMA_signal_3803, n3995}) ) ;
    xnor_HPC2 U4254 ( .a ({new_AGEMA_signal_3492, n4133}), .b ({new_AGEMA_signal_3803, n3995}), .c ({new_AGEMA_signal_4117, n4038}) ) ;
    xnor_HPC2 U4255 ( .a ({new_AGEMA_signal_4117, n4038}), .b ({new_AGEMA_signal_4093, n3996}), .c ({new_AGEMA_signal_4404, n3997}) ) ;
    xnor_HPC2 U4256 ( .a ({new_AGEMA_signal_4404, n3997}), .b ({new_AGEMA_signal_4110, n4027}), .c ({state_out_s1[230], state_out_s0[230]}) ) ;
    xnor_HPC2 U4258 ( .a ({new_AGEMA_signal_4096, n3998}), .b ({new_AGEMA_signal_4111, n4029}), .c ({new_AGEMA_signal_4405, n4000}) ) ;
    xor_HPC2 U4259 ( .a ({new_AGEMA_signal_2797, n3251}), .b ({new_AGEMA_signal_3189, z2[48]}), .c ({new_AGEMA_signal_3493, n4131}) ) ;
    xor_HPC2 U4260 ( .a ({new_AGEMA_signal_3561, z3[48]}), .b ({state_in_s1[200], state_in_s0[200]}), .c ({new_AGEMA_signal_3804, n3999}) ) ;
    xnor_HPC2 U4261 ( .a ({new_AGEMA_signal_3493, n4131}), .b ({new_AGEMA_signal_3804, n3999}), .c ({new_AGEMA_signal_4118, n4058}) ) ;
    xnor_HPC2 U4262 ( .a ({new_AGEMA_signal_4405, n4000}), .b ({new_AGEMA_signal_4118, n4058}), .c ({state_out_s1[231], state_out_s0[231]}) ) ;
    xor_HPC2 U4264 ( .a ({new_AGEMA_signal_2800, n3250}), .b ({new_AGEMA_signal_3196, z2[49]}), .c ({new_AGEMA_signal_3494, n4128}) ) ;
    xor_HPC2 U4265 ( .a ({new_AGEMA_signal_3562, z3[49]}), .b ({state_in_s1[201], state_in_s0[201]}), .c ({new_AGEMA_signal_3805, n4001}) ) ;
    xnor_HPC2 U4266 ( .a ({new_AGEMA_signal_3494, n4128}), .b ({new_AGEMA_signal_3805, n4001}), .c ({new_AGEMA_signal_4119, n4074}) ) ;
    xor_HPC2 U4267 ( .a ({new_AGEMA_signal_4099, n4002}), .b ({new_AGEMA_signal_4112, n4032}), .c ({new_AGEMA_signal_4406, n4003}) ) ;
    xnor_HPC2 U4268 ( .a ({new_AGEMA_signal_4119, n4074}), .b ({new_AGEMA_signal_4406, n4003}), .c ({state_out_s1[216], state_out_s0[216]}) ) ;
    xor_HPC2 U4270 ( .a ({new_AGEMA_signal_2803, n3249}), .b ({new_AGEMA_signal_3195, z2[50]}), .c ({new_AGEMA_signal_3495, n4126}) ) ;
    xnor_HPC2 U4271 ( .a ({new_AGEMA_signal_3564, z3[50]}), .b ({state_in_s1[202], state_in_s0[202]}), .c ({new_AGEMA_signal_3806, n4004}) ) ;
    xnor_HPC2 U4272 ( .a ({new_AGEMA_signal_3495, n4126}), .b ({new_AGEMA_signal_3806, n4004}), .c ({new_AGEMA_signal_4120, n4267}) ) ;
    xor_HPC2 U4273 ( .a ({new_AGEMA_signal_4120, n4267}), .b ({new_AGEMA_signal_4113, n4035}), .c ({new_AGEMA_signal_4407, n4005}) ) ;
    xnor_HPC2 U4274 ( .a ({new_AGEMA_signal_4101, n4006}), .b ({new_AGEMA_signal_4407, n4005}), .c ({state_out_s1[217], state_out_s0[217]}) ) ;
    xnor_HPC2 U4276 ( .a ({new_AGEMA_signal_4114, n4046}), .b ({new_AGEMA_signal_4103, n4007}), .c ({new_AGEMA_signal_4408, n4009}) ) ;
    xor_HPC2 U4277 ( .a ({new_AGEMA_signal_2805, n3248}), .b ({new_AGEMA_signal_3194, z2[51]}), .c ({new_AGEMA_signal_3496, n4125}) ) ;
    xor_HPC2 U4278 ( .a ({new_AGEMA_signal_3565, z3[51]}), .b ({state_in_s1[203], state_in_s0[203]}), .c ({new_AGEMA_signal_3807, n4008}) ) ;
    xnor_HPC2 U4279 ( .a ({new_AGEMA_signal_3496, n4125}), .b ({new_AGEMA_signal_3807, n4008}), .c ({new_AGEMA_signal_4121, n4251}) ) ;
    xnor_HPC2 U4280 ( .a ({new_AGEMA_signal_4408, n4009}), .b ({new_AGEMA_signal_4121, n4251}), .c ({state_out_s1[218], state_out_s0[218]}) ) ;
    xnor_HPC2 U4282 ( .a ({new_AGEMA_signal_4105, n4010}), .b ({new_AGEMA_signal_4115, n4050}), .c ({new_AGEMA_signal_4409, n4012}) ) ;
    xor_HPC2 U4283 ( .a ({new_AGEMA_signal_2807, n3247}), .b ({new_AGEMA_signal_3192, z2[52]}), .c ({new_AGEMA_signal_3497, n4123}) ) ;
    xnor_HPC2 U4284 ( .a ({new_AGEMA_signal_3566, z3[52]}), .b ({state_in_s1[204], state_in_s0[204]}), .c ({new_AGEMA_signal_3808, n4011}) ) ;
    xnor_HPC2 U4285 ( .a ({new_AGEMA_signal_3497, n4123}), .b ({new_AGEMA_signal_3808, n4011}), .c ({new_AGEMA_signal_4122, n4243}) ) ;
    xnor_HPC2 U4286 ( .a ({new_AGEMA_signal_4409, n4012}), .b ({new_AGEMA_signal_4122, n4243}), .c ({state_out_s1[219], state_out_s0[219]}) ) ;
    xor_HPC2 U4288 ( .a ({new_AGEMA_signal_2810, n3246}), .b ({new_AGEMA_signal_3190, z2[53]}), .c ({new_AGEMA_signal_3498, n4120}) ) ;
    xnor_HPC2 U4289 ( .a ({new_AGEMA_signal_3567, z3[53]}), .b ({state_in_s1[205], state_in_s0[205]}), .c ({new_AGEMA_signal_3809, n4013}) ) ;
    xnor_HPC2 U4290 ( .a ({new_AGEMA_signal_3498, n4120}), .b ({new_AGEMA_signal_3809, n4013}), .c ({new_AGEMA_signal_4123, n4233}) ) ;
    xor_HPC2 U4291 ( .a ({new_AGEMA_signal_4123, n4233}), .b ({new_AGEMA_signal_4116, n4055}), .c ({new_AGEMA_signal_4410, n4014}) ) ;
    xnor_HPC2 U4292 ( .a ({new_AGEMA_signal_4106, n4015}), .b ({new_AGEMA_signal_4410, n4014}), .c ({state_out_s1[220], state_out_s0[220]}) ) ;
    xor_HPC2 U4294 ( .a ({new_AGEMA_signal_2813, n3245}), .b ({new_AGEMA_signal_3200, z2[54]}), .c ({new_AGEMA_signal_3499, n4118}) ) ;
    xnor_HPC2 U4295 ( .a ({new_AGEMA_signal_3568, z3[54]}), .b ({state_in_s1[206], state_in_s0[206]}), .c ({new_AGEMA_signal_3810, n4016}) ) ;
    xnor_HPC2 U4296 ( .a ({new_AGEMA_signal_3499, n4118}), .b ({new_AGEMA_signal_3810, n4016}), .c ({new_AGEMA_signal_4124, n4091}) ) ;
    xor_HPC2 U4297 ( .a ({new_AGEMA_signal_4124, n4091}), .b ({new_AGEMA_signal_4117, n4038}), .c ({new_AGEMA_signal_4411, n4017}) ) ;
    xnor_HPC2 U4298 ( .a ({new_AGEMA_signal_4107, n4018}), .b ({new_AGEMA_signal_4411, n4017}), .c ({state_out_s1[221], state_out_s0[221]}) ) ;
    xnor_HPC2 U4300 ( .a ({new_AGEMA_signal_4108, n4019}), .b ({new_AGEMA_signal_4118, n4058}), .c ({new_AGEMA_signal_4412, n4021}) ) ;
    xor_HPC2 U4301 ( .a ({new_AGEMA_signal_2816, n3244}), .b ({new_AGEMA_signal_3197, z2[55]}), .c ({new_AGEMA_signal_3500, n4117}) ) ;
    xor_HPC2 U4302 ( .a ({new_AGEMA_signal_3569, z3[55]}), .b ({state_in_s1[207], state_in_s0[207]}), .c ({new_AGEMA_signal_3811, n4020}) ) ;
    xnor_HPC2 U4303 ( .a ({new_AGEMA_signal_3500, n4117}), .b ({new_AGEMA_signal_3811, n4020}), .c ({new_AGEMA_signal_4125, n4060}) ) ;
    xnor_HPC2 U4304 ( .a ({new_AGEMA_signal_4412, n4021}), .b ({new_AGEMA_signal_4125, n4060}), .c ({state_out_s1[222], state_out_s0[222]}) ) ;
    xor_HPC2 U4306 ( .a ({new_AGEMA_signal_2819, n3243}), .b ({new_AGEMA_signal_3199, z2[56]}), .c ({new_AGEMA_signal_3501, n4114}) ) ;
    xor_HPC2 U4307 ( .a ({new_AGEMA_signal_3570, z3[56]}), .b ({state_in_s1[192], state_in_s0[192]}), .c ({new_AGEMA_signal_3812, n4022}) ) ;
    xnor_HPC2 U4308 ( .a ({new_AGEMA_signal_3501, n4114}), .b ({new_AGEMA_signal_3812, n4022}), .c ({new_AGEMA_signal_4126, n4071}) ) ;
    xnor_HPC2 U4309 ( .a ({new_AGEMA_signal_4109, n4023}), .b ({new_AGEMA_signal_4126, n4071}), .c ({new_AGEMA_signal_4413, n4024}) ) ;
    xnor_HPC2 U4310 ( .a ({new_AGEMA_signal_4413, n4024}), .b ({new_AGEMA_signal_4119, n4074}), .c ({state_out_s1[223], state_out_s0[223]}) ) ;
    xor_HPC2 U4312 ( .a ({new_AGEMA_signal_2821, n3242}), .b ({new_AGEMA_signal_3204, z2[57]}), .c ({new_AGEMA_signal_3502, n4112}) ) ;
    xnor_HPC2 U4313 ( .a ({new_AGEMA_signal_3571, z3[57]}), .b ({state_in_s1[193], state_in_s0[193]}), .c ({new_AGEMA_signal_3813, n4025}) ) ;
    xnor_HPC2 U4314 ( .a ({new_AGEMA_signal_3502, n4112}), .b ({new_AGEMA_signal_3813, n4025}), .c ({new_AGEMA_signal_4127, n4270}) ) ;
    xor_HPC2 U4315 ( .a ({new_AGEMA_signal_4120, n4267}), .b ({new_AGEMA_signal_4127, n4270}), .c ({new_AGEMA_signal_4414, n4026}) ) ;
    xnor_HPC2 U4316 ( .a ({new_AGEMA_signal_4110, n4027}), .b ({new_AGEMA_signal_4414, n4026}), .c ({state_out_s1[208], state_out_s0[208]}) ) ;
    xor_HPC2 U4318 ( .a ({new_AGEMA_signal_2823, n3241}), .b ({new_AGEMA_signal_3203, z2[58]}), .c ({new_AGEMA_signal_3503, n4226}) ) ;
    xnor_HPC2 U4319 ( .a ({new_AGEMA_signal_3572, z3[58]}), .b ({state_in_s1[194], state_in_s0[194]}), .c ({new_AGEMA_signal_3814, n4028}) ) ;
    xnor_HPC2 U4320 ( .a ({new_AGEMA_signal_3503, n4226}), .b ({new_AGEMA_signal_3814, n4028}), .c ({new_AGEMA_signal_4128, n4257}) ) ;
    xnor_HPC2 U4321 ( .a ({new_AGEMA_signal_4128, n4257}), .b ({new_AGEMA_signal_4111, n4029}), .c ({new_AGEMA_signal_4415, n4030}) ) ;
    xnor_HPC2 U4322 ( .a ({new_AGEMA_signal_4415, n4030}), .b ({new_AGEMA_signal_4121, n4251}), .c ({state_out_s1[209], state_out_s0[209]}) ) ;
    xor_HPC2 U4324 ( .a ({new_AGEMA_signal_2825, n3240}), .b ({new_AGEMA_signal_3202, z2[59]}), .c ({new_AGEMA_signal_3504, n4223}) ) ;
    xnor_HPC2 U4325 ( .a ({new_AGEMA_signal_3573, z3[59]}), .b ({state_in_s1[195], state_in_s0[195]}), .c ({new_AGEMA_signal_3815, n4031}) ) ;
    xnor_HPC2 U4326 ( .a ({new_AGEMA_signal_3504, n4223}), .b ({new_AGEMA_signal_3815, n4031}), .c ({new_AGEMA_signal_4129, n4246}) ) ;
    xnor_HPC2 U4327 ( .a ({new_AGEMA_signal_4129, n4246}), .b ({new_AGEMA_signal_4112, n4032}), .c ({new_AGEMA_signal_4416, n4033}) ) ;
    xnor_HPC2 U4328 ( .a ({new_AGEMA_signal_4416, n4033}), .b ({new_AGEMA_signal_4122, n4243}), .c ({state_out_s1[210], state_out_s0[210]}) ) ;
    xor_HPC2 U4330 ( .a ({new_AGEMA_signal_2828, n3238}), .b ({new_AGEMA_signal_3201, z2[60]}), .c ({new_AGEMA_signal_3505, n4220}) ) ;
    xor_HPC2 U4331 ( .a ({new_AGEMA_signal_3575, z3[60]}), .b ({state_in_s1[196], state_in_s0[196]}), .c ({new_AGEMA_signal_3816, n4034}) ) ;
    xnor_HPC2 U4332 ( .a ({new_AGEMA_signal_3505, n4220}), .b ({new_AGEMA_signal_3816, n4034}), .c ({new_AGEMA_signal_4130, n4266}) ) ;
    xor_HPC2 U4333 ( .a ({new_AGEMA_signal_4123, n4233}), .b ({new_AGEMA_signal_4113, n4035}), .c ({new_AGEMA_signal_4417, n4036}) ) ;
    xnor_HPC2 U4334 ( .a ({new_AGEMA_signal_4130, n4266}), .b ({new_AGEMA_signal_4417, n4036}), .c ({state_out_s1[211], state_out_s0[211]}) ) ;
    xnor_HPC2 U4336 ( .a ({new_AGEMA_signal_3206, z2[0]}), .b ({new_AGEMA_signal_2831, n4041}), .c ({new_AGEMA_signal_3506, n4099}) ) ;
    xnor_HPC2 U4337 ( .a ({1'b0, rcon[0]}), .b ({new_AGEMA_signal_3506, n4099}), .c ({new_AGEMA_signal_3817, n4224}) ) ;
    xnor_HPC2 U4338 ( .a ({new_AGEMA_signal_3817, n4224}), .b ({new_AGEMA_signal_3519, z3[0]}), .c ({new_AGEMA_signal_4131, n4037}) ) ;
    xnor_HPC2 U4339 ( .a ({new_AGEMA_signal_4131, n4037}), .b ({state_in_s1[248], state_in_s0[248]}), .c ({new_AGEMA_signal_4418, n4092}) ) ;
    xnor_HPC2 U4340 ( .a ({new_AGEMA_signal_4418, n4092}), .b ({new_AGEMA_signal_4127, n4270}), .c ({new_AGEMA_signal_4550, n4039}) ) ;
    xnor_HPC2 U4341 ( .a ({new_AGEMA_signal_4550, n4039}), .b ({new_AGEMA_signal_4117, n4038}), .c ({state_out_s1[215], state_out_s0[215]}) ) ;
    xor_HPC2 U4342 ( .a ({new_AGEMA_signal_4418, n4092}), .b ({new_AGEMA_signal_4102, n4095}), .c ({new_AGEMA_signal_4551, n4040}) ) ;
    xnor_HPC2 U4343 ( .a ({new_AGEMA_signal_4083, n4269}), .b ({new_AGEMA_signal_4551, n4040}), .c ({state_out_s1[248], state_out_s0[248]}) ) ;
    xnor_HPC2 U4347 ( .a ({new_AGEMA_signal_2834, n3237}), .b ({new_AGEMA_signal_3294, z2[8]}), .c ({new_AGEMA_signal_3507, n4202}) ) ;
    xor_HPC2 U4348 ( .a ({new_AGEMA_signal_3581, z3[8]}), .b ({state_in_s1[240], state_in_s0[240]}), .c ({new_AGEMA_signal_3818, n4042}) ) ;
    xnor_HPC2 U4349 ( .a ({new_AGEMA_signal_3507, n4202}), .b ({new_AGEMA_signal_3818, n4042}), .c ({new_AGEMA_signal_4132, n4061}) ) ;
    xnor_HPC2 U4350 ( .a ({new_AGEMA_signal_4104, n4063}), .b ({new_AGEMA_signal_4132, n4061}), .c ({new_AGEMA_signal_4419, n4043}) ) ;
    xnor_HPC2 U4351 ( .a ({new_AGEMA_signal_4098, n4044}), .b ({new_AGEMA_signal_4419, n4043}), .c ({state_out_s1[240], state_out_s0[240]}) ) ;
    xor_HPC2 U4353 ( .a ({new_AGEMA_signal_2837, n3236}), .b ({new_AGEMA_signal_3198, z2[61]}), .c ({new_AGEMA_signal_3508, n4215}) ) ;
    xnor_HPC2 U4354 ( .a ({new_AGEMA_signal_3576, z3[61]}), .b ({state_in_s1[197], state_in_s0[197]}), .c ({new_AGEMA_signal_3819, n4045}) ) ;
    xnor_HPC2 U4355 ( .a ({new_AGEMA_signal_3508, n4215}), .b ({new_AGEMA_signal_3819, n4045}), .c ({new_AGEMA_signal_4133, n4253}) ) ;
    xnor_HPC2 U4356 ( .a ({new_AGEMA_signal_4133, n4253}), .b ({new_AGEMA_signal_4124, n4091}), .c ({new_AGEMA_signal_4420, n4047}) ) ;
    xnor_HPC2 U4357 ( .a ({new_AGEMA_signal_4420, n4047}), .b ({new_AGEMA_signal_4114, n4046}), .c ({state_out_s1[212], state_out_s0[212]}) ) ;
    xor_HPC2 U4359 ( .a ({new_AGEMA_signal_2840, n3235}), .b ({new_AGEMA_signal_3209, z2[62]}), .c ({new_AGEMA_signal_3509, n4107}) ) ;
    xnor_HPC2 U4360 ( .a ({new_AGEMA_signal_3509, n4107}), .b ({new_AGEMA_signal_3577, z3[62]}), .c ({new_AGEMA_signal_3820, n4048}) ) ;
    xnor_HPC2 U4361 ( .a ({new_AGEMA_signal_3820, n4048}), .b ({state_in_s1[198], state_in_s0[198]}), .c ({new_AGEMA_signal_4134, n4242}) ) ;
    xnor_HPC2 U4362 ( .a ({new_AGEMA_signal_4132, n4061}), .b ({new_AGEMA_signal_4134, n4242}), .c ({new_AGEMA_signal_4421, n4049}) ) ;
    xnor_HPC2 U4363 ( .a ({new_AGEMA_signal_4097, n4239}), .b ({new_AGEMA_signal_4421, n4049}), .c ({state_out_s1[198], state_out_s0[198]}) ) ;
    xor_HPC2 U4364 ( .a ({new_AGEMA_signal_4115, n4050}), .b ({new_AGEMA_signal_4134, n4242}), .c ({new_AGEMA_signal_4422, n4051}) ) ;
    xnor_HPC2 U4365 ( .a ({new_AGEMA_signal_4125, n4060}), .b ({new_AGEMA_signal_4422, n4051}), .c ({state_out_s1[213], state_out_s0[213]}) ) ;
    xor_HPC2 U4369 ( .a ({new_AGEMA_signal_3208, z2[4]}), .b ({new_AGEMA_signal_2990, n3232}), .c ({new_AGEMA_signal_3510, n4250}) ) ;
    xor_HPC2 U4370 ( .a ({new_AGEMA_signal_2846, n3234}), .b ({new_AGEMA_signal_3205, z2[63]}), .c ({new_AGEMA_signal_3511, n4104}) ) ;
    xor_HPC2 U4371 ( .a ({new_AGEMA_signal_3511, n4104}), .b ({new_AGEMA_signal_3509, n4107}), .c ({new_AGEMA_signal_3821, n4052}) ) ;
    xnor_HPC2 U4372 ( .a ({new_AGEMA_signal_3510, n4250}), .b ({new_AGEMA_signal_3821, n4052}), .c ({state_out_s1[134], state_out_s0[134]}) ) ;
    xnor_HPC2 U4373 ( .a ({new_AGEMA_signal_4079, n4072}), .b ({new_AGEMA_signal_4100, n4229}), .c ({new_AGEMA_signal_4423, n4054}) ) ;
    xnor_HPC2 U4374 ( .a ({new_AGEMA_signal_3578, z3[63]}), .b ({state_in_s1[199], state_in_s0[199]}), .c ({new_AGEMA_signal_3822, n4053}) ) ;
    xnor_HPC2 U4375 ( .a ({new_AGEMA_signal_3511, n4104}), .b ({new_AGEMA_signal_3822, n4053}), .c ({new_AGEMA_signal_4136, n4232}) ) ;
    xnor_HPC2 U4376 ( .a ({new_AGEMA_signal_4423, n4054}), .b ({new_AGEMA_signal_4136, n4232}), .c ({state_out_s1[199], state_out_s0[199]}) ) ;
    xor_HPC2 U4377 ( .a ({new_AGEMA_signal_4136, n4232}), .b ({new_AGEMA_signal_4116, n4055}), .c ({new_AGEMA_signal_4424, n4056}) ) ;
    xnor_HPC2 U4378 ( .a ({new_AGEMA_signal_4126, n4071}), .b ({new_AGEMA_signal_4424, n4056}), .c ({state_out_s1[214], state_out_s0[214]}) ) ;
    xnor_HPC2 U4382 ( .a ({new_AGEMA_signal_3212, z2[1]}), .b ({new_AGEMA_signal_2849, n4066}), .c ({new_AGEMA_signal_3512, n4101}) ) ;
    xnor_HPC2 U4383 ( .a ({1'b0, n4206}), .b ({new_AGEMA_signal_3512, n4101}), .c ({new_AGEMA_signal_3823, n4222}) ) ;
    xor_HPC2 U4384 ( .a ({new_AGEMA_signal_3823, n4222}), .b ({new_AGEMA_signal_3530, z3[1]}), .c ({new_AGEMA_signal_4137, n4057}) ) ;
    xnor_HPC2 U4385 ( .a ({state_in_s1[249], state_in_s0[249]}), .b ({new_AGEMA_signal_4137, n4057}), .c ({new_AGEMA_signal_4425, n4065}) ) ;
    xnor_HPC2 U4386 ( .a ({new_AGEMA_signal_4128, n4257}), .b ({new_AGEMA_signal_4425, n4065}), .c ({new_AGEMA_signal_4558, n4059}) ) ;
    xnor_HPC2 U4387 ( .a ({new_AGEMA_signal_4558, n4059}), .b ({new_AGEMA_signal_4118, n4058}), .c ({state_out_s1[200], state_out_s0[200]}) ) ;
    xnor_HPC2 U4388 ( .a ({new_AGEMA_signal_4132, n4061}), .b ({new_AGEMA_signal_4125, n4060}), .c ({new_AGEMA_signal_4426, n4062}) ) ;
    xnor_HPC2 U4389 ( .a ({new_AGEMA_signal_4426, n4062}), .b ({new_AGEMA_signal_4425, n4065}), .c ({state_out_s1[207], state_out_s0[207]}) ) ;
    xor_HPC2 U4390 ( .a ({new_AGEMA_signal_4085, n4258}), .b ({new_AGEMA_signal_4104, n4063}), .c ({new_AGEMA_signal_4427, n4064}) ) ;
    xnor_HPC2 U4391 ( .a ({new_AGEMA_signal_4425, n4065}), .b ({new_AGEMA_signal_4427, n4064}), .c ({state_out_s1[249], state_out_s0[249]}) ) ;
    xnor_HPC2 U4397 ( .a ({new_AGEMA_signal_3211, z2[2]}), .b ({new_AGEMA_signal_3824, n3287}), .c ({new_AGEMA_signal_4138, n4217}) ) ;
    xnor_HPC2 U4398 ( .a ({new_AGEMA_signal_3541, z3[2]}), .b ({state_in_s1[250], state_in_s0[250]}), .c ({new_AGEMA_signal_3825, n4070}) ) ;
    xnor_HPC2 U4399 ( .a ({new_AGEMA_signal_4138, n4217}), .b ({new_AGEMA_signal_3825, n4070}), .c ({new_AGEMA_signal_4428, n4078}) ) ;
    xnor_HPC2 U4400 ( .a ({new_AGEMA_signal_4079, n4072}), .b ({new_AGEMA_signal_4126, n4071}), .c ({new_AGEMA_signal_4429, n4073}) ) ;
    xnor_HPC2 U4401 ( .a ({new_AGEMA_signal_4428, n4078}), .b ({new_AGEMA_signal_4429, n4073}), .c ({state_out_s1[192], state_out_s0[192]}) ) ;
    xnor_HPC2 U4402 ( .a ({new_AGEMA_signal_4129, n4246}), .b ({new_AGEMA_signal_4119, n4074}), .c ({new_AGEMA_signal_4430, n4075}) ) ;
    xnor_HPC2 U4403 ( .a ({new_AGEMA_signal_4428, n4078}), .b ({new_AGEMA_signal_4430, n4075}), .c ({state_out_s1[201], state_out_s0[201]}) ) ;
    xnor_HPC2 U4404 ( .a ({new_AGEMA_signal_4088, n4245}), .b ({new_AGEMA_signal_4080, n4076}), .c ({new_AGEMA_signal_4431, n4077}) ) ;
    xnor_HPC2 U4405 ( .a ({new_AGEMA_signal_4428, n4078}), .b ({new_AGEMA_signal_4431, n4077}), .c ({state_out_s1[250], state_out_s0[250]}) ) ;
    xnor_HPC2 U4410 ( .a ({new_AGEMA_signal_3210, z2[3]}), .b ({new_AGEMA_signal_4432, n3233}), .c ({new_AGEMA_signal_4564, n4262}) ) ;
    xnor_HPC2 U4411 ( .a ({new_AGEMA_signal_3508, n4215}), .b ({new_AGEMA_signal_4564, n4262}), .c ({new_AGEMA_signal_4602, n4082}) ) ;
    xnor_HPC2 U4412 ( .a ({new_AGEMA_signal_4602, n4082}), .b ({new_AGEMA_signal_3509, n4107}), .c ({state_out_s1[133], state_out_s0[133]}) ) ;
    xnor_HPC2 U4413 ( .a ({new_AGEMA_signal_4564, n4262}), .b ({new_AGEMA_signal_4138, n4217}), .c ({new_AGEMA_signal_4603, n4083}) ) ;
    xnor_HPC2 U4414 ( .a ({new_AGEMA_signal_4603, n4083}), .b ({new_AGEMA_signal_3507, n4202}), .c ({state_out_s1[186], state_out_s0[186]}) ) ;
    xor_HPC2 U4419 ( .a ({new_AGEMA_signal_4433, n3239}), .b ({new_AGEMA_signal_3269, z2[7]}), .c ({new_AGEMA_signal_4565, n4219}) ) ;
    xnor_HPC2 U4420 ( .a ({new_AGEMA_signal_4565, n4219}), .b ({new_AGEMA_signal_3463, n4192}), .c ({new_AGEMA_signal_4604, n4088}) ) ;
    xnor_HPC2 U4421 ( .a ({new_AGEMA_signal_3826, n3230}), .b ({new_AGEMA_signal_3272, z2[6]}), .c ({new_AGEMA_signal_4143, n4228}) ) ;
    xnor_HPC2 U4422 ( .a ({new_AGEMA_signal_4604, n4088}), .b ({new_AGEMA_signal_4143, n4228}), .c ({state_out_s1[190], state_out_s0[190]}) ) ;
    xnor_HPC2 U4423 ( .a ({new_AGEMA_signal_3580, z3[7]}), .b ({state_in_s1[255], state_in_s0[255]}), .c ({new_AGEMA_signal_3827, n4089}) ) ;
    xnor_HPC2 U4424 ( .a ({new_AGEMA_signal_4565, n4219}), .b ({new_AGEMA_signal_3827, n4089}), .c ({new_AGEMA_signal_4605, n4097}) ) ;
    xnor_HPC2 U4425 ( .a ({new_AGEMA_signal_4133, n4253}), .b ({new_AGEMA_signal_4605, n4097}), .c ({new_AGEMA_signal_4627, n4090}) ) ;
    xnor_HPC2 U4426 ( .a ({new_AGEMA_signal_4094, n4255}), .b ({new_AGEMA_signal_4627, n4090}), .c ({state_out_s1[197], state_out_s0[197]}) ) ;
    xnor_HPC2 U4427 ( .a ({new_AGEMA_signal_4605, n4097}), .b ({new_AGEMA_signal_4124, n4091}), .c ({new_AGEMA_signal_4628, n4093}) ) ;
    xnor_HPC2 U4428 ( .a ({new_AGEMA_signal_4628, n4093}), .b ({new_AGEMA_signal_4418, n4092}), .c ({state_out_s1[206], state_out_s0[206]}) ) ;
    xnor_HPC2 U4429 ( .a ({new_AGEMA_signal_4102, n4095}), .b ({new_AGEMA_signal_4095, n4094}), .c ({new_AGEMA_signal_4434, n4096}) ) ;
    xnor_HPC2 U4430 ( .a ({new_AGEMA_signal_4605, n4097}), .b ({new_AGEMA_signal_4434, n4096}), .c ({state_out_s1[255], state_out_s0[255]}) ) ;
    xnor_HPC2 U4431 ( .a ({new_AGEMA_signal_3511, n4104}), .b ({new_AGEMA_signal_3506, n4099}), .c ({new_AGEMA_signal_3828, n4098}) ) ;
    xnor_HPC2 U4433 ( .a ({new_AGEMA_signal_3207, z2[5]}), .b ({new_AGEMA_signal_2858, n4103}), .c ({new_AGEMA_signal_3514, n4205}) ) ;
    xnor_HPC2 U4434 ( .a ({1'b0, rcon[1]}), .b ({new_AGEMA_signal_3514, n4205}), .c ({new_AGEMA_signal_3829, n4210}) ) ;
    xnor_HPC2 U4435 ( .a ({new_AGEMA_signal_3828, n4098}), .b ({new_AGEMA_signal_3829, n4210}), .c ({state_out_s1[135], state_out_s0[135]}) ) ;
    xor_HPC2 U4436 ( .a ({new_AGEMA_signal_3506, n4099}), .b ({new_AGEMA_signal_4143, n4228}), .c ({new_AGEMA_signal_4435, n4100}) ) ;
    xnor_HPC2 U4437 ( .a ({new_AGEMA_signal_3512, n4101}), .b ({new_AGEMA_signal_4435, n4100}), .c ({new_AGEMA_signal_4566, n4102}) ) ;
    xnor_HPC2 U4438 ( .a ({1'b0, rcon[1]}), .b ({new_AGEMA_signal_4566, n4102}), .c ({state_out_s1[184], state_out_s0[184]}) ) ;
    xor_HPC2 U4440 ( .a ({new_AGEMA_signal_3502, n4112}), .b ({new_AGEMA_signal_3511, n4104}), .c ({new_AGEMA_signal_3830, n4105}) ) ;
    xnor_HPC2 U4441 ( .a ({new_AGEMA_signal_3503, n4226}), .b ({new_AGEMA_signal_3830, n4105}), .c ({state_out_s1[129], state_out_s0[129]}) ) ;
    xor_HPC2 U4442 ( .a ({new_AGEMA_signal_3502, n4112}), .b ({new_AGEMA_signal_3501, n4114}), .c ({new_AGEMA_signal_3831, n4106}) ) ;
    xnor_HPC2 U4443 ( .a ({new_AGEMA_signal_3509, n4107}), .b ({new_AGEMA_signal_3831, n4106}), .c ({state_out_s1[128], state_out_s0[128]}) ) ;
    xor_HPC2 U4444 ( .a ({new_AGEMA_signal_3508, n4215}), .b ({new_AGEMA_signal_3501, n4114}), .c ({new_AGEMA_signal_3832, n4108}) ) ;
    xnor_HPC2 U4445 ( .a ({new_AGEMA_signal_3500, n4117}), .b ({new_AGEMA_signal_3832, n4108}), .c ({state_out_s1[143], state_out_s0[143]}) ) ;
    xor_HPC2 U4446 ( .a ({new_AGEMA_signal_3499, n4118}), .b ({new_AGEMA_signal_3505, n4220}), .c ({new_AGEMA_signal_3833, n4109}) ) ;
    xnor_HPC2 U4447 ( .a ({new_AGEMA_signal_3500, n4117}), .b ({new_AGEMA_signal_3833, n4109}), .c ({state_out_s1[142], state_out_s0[142]}) ) ;
    xor_HPC2 U4448 ( .a ({new_AGEMA_signal_3499, n4118}), .b ({new_AGEMA_signal_3504, n4223}), .c ({new_AGEMA_signal_3834, n4110}) ) ;
    xnor_HPC2 U4449 ( .a ({new_AGEMA_signal_3498, n4120}), .b ({new_AGEMA_signal_3834, n4110}), .c ({state_out_s1[141], state_out_s0[141]}) ) ;
    xor_HPC2 U4450 ( .a ({new_AGEMA_signal_3498, n4120}), .b ({new_AGEMA_signal_3497, n4123}), .c ({new_AGEMA_signal_3835, n4111}) ) ;
    xnor_HPC2 U4451 ( .a ({new_AGEMA_signal_3503, n4226}), .b ({new_AGEMA_signal_3835, n4111}), .c ({state_out_s1[140], state_out_s0[140]}) ) ;
    xor_HPC2 U4452 ( .a ({new_AGEMA_signal_3502, n4112}), .b ({new_AGEMA_signal_3496, n4125}), .c ({new_AGEMA_signal_3836, n4113}) ) ;
    xnor_HPC2 U4453 ( .a ({new_AGEMA_signal_3497, n4123}), .b ({new_AGEMA_signal_3836, n4113}), .c ({state_out_s1[139], state_out_s0[139]}) ) ;
    xor_HPC2 U4454 ( .a ({new_AGEMA_signal_3495, n4126}), .b ({new_AGEMA_signal_3501, n4114}), .c ({new_AGEMA_signal_3837, n4115}) ) ;
    xnor_HPC2 U4455 ( .a ({new_AGEMA_signal_3496, n4125}), .b ({new_AGEMA_signal_3837, n4115}), .c ({state_out_s1[138], state_out_s0[138]}) ) ;
    xor_HPC2 U4456 ( .a ({new_AGEMA_signal_3495, n4126}), .b ({new_AGEMA_signal_3494, n4128}), .c ({new_AGEMA_signal_3838, n4116}) ) ;
    xnor_HPC2 U4457 ( .a ({new_AGEMA_signal_3500, n4117}), .b ({new_AGEMA_signal_3838, n4116}), .c ({state_out_s1[137], state_out_s0[137]}) ) ;
    xor_HPC2 U4458 ( .a ({new_AGEMA_signal_3499, n4118}), .b ({new_AGEMA_signal_3494, n4128}), .c ({new_AGEMA_signal_3839, n4119}) ) ;
    xnor_HPC2 U4459 ( .a ({new_AGEMA_signal_3493, n4131}), .b ({new_AGEMA_signal_3839, n4119}), .c ({state_out_s1[136], state_out_s0[136]}) ) ;
    xor_HPC2 U4460 ( .a ({new_AGEMA_signal_3498, n4120}), .b ({new_AGEMA_signal_3492, n4133}), .c ({new_AGEMA_signal_3840, n4121}) ) ;
    xnor_HPC2 U4461 ( .a ({new_AGEMA_signal_3493, n4131}), .b ({new_AGEMA_signal_3840, n4121}), .c ({state_out_s1[151], state_out_s0[151]}) ) ;
    xor_HPC2 U4462 ( .a ({new_AGEMA_signal_3491, n4135}), .b ({new_AGEMA_signal_3492, n4133}), .c ({new_AGEMA_signal_3841, n4122}) ) ;
    xnor_HPC2 U4463 ( .a ({new_AGEMA_signal_3497, n4123}), .b ({new_AGEMA_signal_3841, n4122}), .c ({state_out_s1[150], state_out_s0[150]}) ) ;
    xor_HPC2 U4464 ( .a ({new_AGEMA_signal_3490, n4137}), .b ({new_AGEMA_signal_3491, n4135}), .c ({new_AGEMA_signal_3842, n4124}) ) ;
    xnor_HPC2 U4465 ( .a ({new_AGEMA_signal_3496, n4125}), .b ({new_AGEMA_signal_3842, n4124}), .c ({state_out_s1[149], state_out_s0[149]}) ) ;
    xor_HPC2 U4466 ( .a ({new_AGEMA_signal_3495, n4126}), .b ({new_AGEMA_signal_3489, n4139}), .c ({new_AGEMA_signal_3843, n4127}) ) ;
    xnor_HPC2 U4467 ( .a ({new_AGEMA_signal_3490, n4137}), .b ({new_AGEMA_signal_3843, n4127}), .c ({state_out_s1[148], state_out_s0[148]}) ) ;
    xor_HPC2 U4468 ( .a ({new_AGEMA_signal_3494, n4128}), .b ({new_AGEMA_signal_3488, n4141}), .c ({new_AGEMA_signal_3844, n4129}) ) ;
    xnor_HPC2 U4469 ( .a ({new_AGEMA_signal_3489, n4139}), .b ({new_AGEMA_signal_3844, n4129}), .c ({state_out_s1[147], state_out_s0[147]}) ) ;
    xor_HPC2 U4470 ( .a ({new_AGEMA_signal_3487, n4143}), .b ({new_AGEMA_signal_3488, n4141}), .c ({new_AGEMA_signal_3845, n4130}) ) ;
    xnor_HPC2 U4471 ( .a ({new_AGEMA_signal_3493, n4131}), .b ({new_AGEMA_signal_3845, n4130}), .c ({state_out_s1[146], state_out_s0[146]}) ) ;
    xor_HPC2 U4472 ( .a ({new_AGEMA_signal_3486, n4145}), .b ({new_AGEMA_signal_3487, n4143}), .c ({new_AGEMA_signal_3846, n4132}) ) ;
    xnor_HPC2 U4473 ( .a ({new_AGEMA_signal_3492, n4133}), .b ({new_AGEMA_signal_3846, n4132}), .c ({state_out_s1[145], state_out_s0[145]}) ) ;
    xor_HPC2 U4474 ( .a ({new_AGEMA_signal_3485, n4147}), .b ({new_AGEMA_signal_3486, n4145}), .c ({new_AGEMA_signal_3847, n4134}) ) ;
    xnor_HPC2 U4475 ( .a ({new_AGEMA_signal_3491, n4135}), .b ({new_AGEMA_signal_3847, n4134}), .c ({state_out_s1[144], state_out_s0[144]}) ) ;
    xor_HPC2 U4476 ( .a ({new_AGEMA_signal_3484, n4149}), .b ({new_AGEMA_signal_3485, n4147}), .c ({new_AGEMA_signal_3848, n4136}) ) ;
    xnor_HPC2 U4477 ( .a ({new_AGEMA_signal_3490, n4137}), .b ({new_AGEMA_signal_3848, n4136}), .c ({state_out_s1[159], state_out_s0[159]}) ) ;
    xor_HPC2 U4478 ( .a ({new_AGEMA_signal_3483, n4151}), .b ({new_AGEMA_signal_3484, n4149}), .c ({new_AGEMA_signal_3849, n4138}) ) ;
    xnor_HPC2 U4479 ( .a ({new_AGEMA_signal_3489, n4139}), .b ({new_AGEMA_signal_3849, n4138}), .c ({state_out_s1[158], state_out_s0[158]}) ) ;
    xor_HPC2 U4480 ( .a ({new_AGEMA_signal_3482, n4153}), .b ({new_AGEMA_signal_3483, n4151}), .c ({new_AGEMA_signal_3850, n4140}) ) ;
    xnor_HPC2 U4481 ( .a ({new_AGEMA_signal_3488, n4141}), .b ({new_AGEMA_signal_3850, n4140}), .c ({state_out_s1[157], state_out_s0[157]}) ) ;
    xor_HPC2 U4482 ( .a ({new_AGEMA_signal_3481, n4155}), .b ({new_AGEMA_signal_3482, n4153}), .c ({new_AGEMA_signal_3851, n4142}) ) ;
    xnor_HPC2 U4483 ( .a ({new_AGEMA_signal_3487, n4143}), .b ({new_AGEMA_signal_3851, n4142}), .c ({state_out_s1[156], state_out_s0[156]}) ) ;
    xor_HPC2 U4484 ( .a ({new_AGEMA_signal_3480, n4157}), .b ({new_AGEMA_signal_3481, n4155}), .c ({new_AGEMA_signal_3852, n4144}) ) ;
    xnor_HPC2 U4485 ( .a ({new_AGEMA_signal_3486, n4145}), .b ({new_AGEMA_signal_3852, n4144}), .c ({state_out_s1[155], state_out_s0[155]}) ) ;
    xor_HPC2 U4486 ( .a ({new_AGEMA_signal_3478, n4159}), .b ({new_AGEMA_signal_3480, n4157}), .c ({new_AGEMA_signal_3853, n4146}) ) ;
    xnor_HPC2 U4487 ( .a ({new_AGEMA_signal_3485, n4147}), .b ({new_AGEMA_signal_3853, n4146}), .c ({state_out_s1[154], state_out_s0[154]}) ) ;
    xor_HPC2 U4488 ( .a ({new_AGEMA_signal_3476, n4161}), .b ({new_AGEMA_signal_3478, n4159}), .c ({new_AGEMA_signal_3854, n4148}) ) ;
    xnor_HPC2 U4489 ( .a ({new_AGEMA_signal_3484, n4149}), .b ({new_AGEMA_signal_3854, n4148}), .c ({state_out_s1[153], state_out_s0[153]}) ) ;
    xor_HPC2 U4490 ( .a ({new_AGEMA_signal_3474, n4163}), .b ({new_AGEMA_signal_3476, n4161}), .c ({new_AGEMA_signal_3855, n4150}) ) ;
    xnor_HPC2 U4491 ( .a ({new_AGEMA_signal_3483, n4151}), .b ({new_AGEMA_signal_3855, n4150}), .c ({state_out_s1[152], state_out_s0[152]}) ) ;
    xor_HPC2 U4492 ( .a ({new_AGEMA_signal_3471, n4164}), .b ({new_AGEMA_signal_3474, n4163}), .c ({new_AGEMA_signal_3856, n4152}) ) ;
    xnor_HPC2 U4493 ( .a ({new_AGEMA_signal_3482, n4153}), .b ({new_AGEMA_signal_3856, n4152}), .c ({state_out_s1[167], state_out_s0[167]}) ) ;
    xor_HPC2 U4494 ( .a ({new_AGEMA_signal_3468, n4166}), .b ({new_AGEMA_signal_3471, n4164}), .c ({new_AGEMA_signal_3857, n4154}) ) ;
    xnor_HPC2 U4495 ( .a ({new_AGEMA_signal_3481, n4155}), .b ({new_AGEMA_signal_3857, n4154}), .c ({state_out_s1[166], state_out_s0[166]}) ) ;
    xor_HPC2 U4496 ( .a ({new_AGEMA_signal_3465, n4169}), .b ({new_AGEMA_signal_3468, n4166}), .c ({new_AGEMA_signal_3858, n4156}) ) ;
    xnor_HPC2 U4497 ( .a ({new_AGEMA_signal_3480, n4157}), .b ({new_AGEMA_signal_3858, n4156}), .c ({state_out_s1[165], state_out_s0[165]}) ) ;
    xor_HPC2 U4498 ( .a ({new_AGEMA_signal_3462, n4170}), .b ({new_AGEMA_signal_3465, n4169}), .c ({new_AGEMA_signal_3859, n4158}) ) ;
    xnor_HPC2 U4499 ( .a ({new_AGEMA_signal_3478, n4159}), .b ({new_AGEMA_signal_3859, n4158}), .c ({state_out_s1[164], state_out_s0[164]}) ) ;
    xor_HPC2 U4500 ( .a ({new_AGEMA_signal_3459, n4172}), .b ({new_AGEMA_signal_3462, n4170}), .c ({new_AGEMA_signal_3860, n4160}) ) ;
    xnor_HPC2 U4501 ( .a ({new_AGEMA_signal_3476, n4161}), .b ({new_AGEMA_signal_3860, n4160}), .c ({state_out_s1[163], state_out_s0[163]}) ) ;
    xor_HPC2 U4502 ( .a ({new_AGEMA_signal_3456, n4174}), .b ({new_AGEMA_signal_3459, n4172}), .c ({new_AGEMA_signal_3861, n4162}) ) ;
    xnor_HPC2 U4503 ( .a ({new_AGEMA_signal_3474, n4163}), .b ({new_AGEMA_signal_3861, n4162}), .c ({state_out_s1[162], state_out_s0[162]}) ) ;
    xor_HPC2 U4504 ( .a ({new_AGEMA_signal_3456, n4174}), .b ({new_AGEMA_signal_3471, n4164}), .c ({new_AGEMA_signal_3862, n4165}) ) ;
    xnor_HPC2 U4505 ( .a ({new_AGEMA_signal_3473, n4177}), .b ({new_AGEMA_signal_3862, n4165}), .c ({state_out_s1[161], state_out_s0[161]}) ) ;
    xor_HPC2 U4506 ( .a ({new_AGEMA_signal_3470, n4178}), .b ({new_AGEMA_signal_3468, n4166}), .c ({new_AGEMA_signal_3863, n4167}) ) ;
    xnor_HPC2 U4507 ( .a ({new_AGEMA_signal_3473, n4177}), .b ({new_AGEMA_signal_3863, n4167}), .c ({state_out_s1[160], state_out_s0[160]}) ) ;
    xor_HPC2 U4508 ( .a ({new_AGEMA_signal_3470, n4178}), .b ({new_AGEMA_signal_3466, n4180}), .c ({new_AGEMA_signal_3864, n4168}) ) ;
    xnor_HPC2 U4509 ( .a ({new_AGEMA_signal_3465, n4169}), .b ({new_AGEMA_signal_3864, n4168}), .c ({state_out_s1[175], state_out_s0[175]}) ) ;
    xor_HPC2 U4510 ( .a ({new_AGEMA_signal_3466, n4180}), .b ({new_AGEMA_signal_3462, n4170}), .c ({new_AGEMA_signal_3865, n4171}) ) ;
    xnor_HPC2 U4511 ( .a ({new_AGEMA_signal_3464, n4183}), .b ({new_AGEMA_signal_3865, n4171}), .c ({state_out_s1[174], state_out_s0[174]}) ) ;
    xor_HPC2 U4512 ( .a ({new_AGEMA_signal_3459, n4172}), .b ({new_AGEMA_signal_3461, n4184}), .c ({new_AGEMA_signal_3866, n4173}) ) ;
    xnor_HPC2 U4513 ( .a ({new_AGEMA_signal_3464, n4183}), .b ({new_AGEMA_signal_3866, n4173}), .c ({state_out_s1[173], state_out_s0[173]}) ) ;
    xor_HPC2 U4514 ( .a ({new_AGEMA_signal_3457, n4186}), .b ({new_AGEMA_signal_3456, n4174}), .c ({new_AGEMA_signal_3867, n4175}) ) ;
    xnor_HPC2 U4515 ( .a ({new_AGEMA_signal_3461, n4184}), .b ({new_AGEMA_signal_3867, n4175}), .c ({state_out_s1[172], state_out_s0[172]}) ) ;
    xor_HPC2 U4516 ( .a ({new_AGEMA_signal_3457, n4186}), .b ({new_AGEMA_signal_3455, n4189}), .c ({new_AGEMA_signal_3868, n4176}) ) ;
    xnor_HPC2 U4517 ( .a ({new_AGEMA_signal_3473, n4177}), .b ({new_AGEMA_signal_3868, n4176}), .c ({state_out_s1[171], state_out_s0[171]}) ) ;
    xor_HPC2 U4518 ( .a ({new_AGEMA_signal_3470, n4178}), .b ({new_AGEMA_signal_3455, n4189}), .c ({new_AGEMA_signal_3869, n4179}) ) ;
    xnor_HPC2 U4519 ( .a ({new_AGEMA_signal_3479, n4191}), .b ({new_AGEMA_signal_3869, n4179}), .c ({state_out_s1[170], state_out_s0[170]}) ) ;
    xor_HPC2 U4520 ( .a ({new_AGEMA_signal_3477, n4193}), .b ({new_AGEMA_signal_3466, n4180}), .c ({new_AGEMA_signal_3870, n4181}) ) ;
    xnor_HPC2 U4521 ( .a ({new_AGEMA_signal_3479, n4191}), .b ({new_AGEMA_signal_3870, n4181}), .c ({state_out_s1[169], state_out_s0[169]}) ) ;
    xor_HPC2 U4522 ( .a ({new_AGEMA_signal_3477, n4193}), .b ({new_AGEMA_signal_3475, n4195}), .c ({new_AGEMA_signal_3871, n4182}) ) ;
    xnor_HPC2 U4523 ( .a ({new_AGEMA_signal_3464, n4183}), .b ({new_AGEMA_signal_3871, n4182}), .c ({state_out_s1[168], state_out_s0[168]}) ) ;
    xor_HPC2 U4524 ( .a ({new_AGEMA_signal_3475, n4195}), .b ({new_AGEMA_signal_3461, n4184}), .c ({new_AGEMA_signal_3872, n4185}) ) ;
    xnor_HPC2 U4525 ( .a ({new_AGEMA_signal_3472, n4198}), .b ({new_AGEMA_signal_3872, n4185}), .c ({state_out_s1[183], state_out_s0[183]}) ) ;
    xor_HPC2 U4526 ( .a ({new_AGEMA_signal_3469, n4199}), .b ({new_AGEMA_signal_3457, n4186}), .c ({new_AGEMA_signal_3873, n4187}) ) ;
    xnor_HPC2 U4527 ( .a ({new_AGEMA_signal_3472, n4198}), .b ({new_AGEMA_signal_3873, n4187}), .c ({state_out_s1[182], state_out_s0[182]}) ) ;
    xor_HPC2 U4528 ( .a ({new_AGEMA_signal_3469, n4199}), .b ({new_AGEMA_signal_3467, n4201}), .c ({new_AGEMA_signal_3874, n4188}) ) ;
    xnor_HPC2 U4529 ( .a ({new_AGEMA_signal_3455, n4189}), .b ({new_AGEMA_signal_3874, n4188}), .c ({state_out_s1[181], state_out_s0[181]}) ) ;
    xor_HPC2 U4530 ( .a ({new_AGEMA_signal_3467, n4201}), .b ({new_AGEMA_signal_3463, n4192}), .c ({new_AGEMA_signal_3875, n4190}) ) ;
    xnor_HPC2 U4531 ( .a ({new_AGEMA_signal_3479, n4191}), .b ({new_AGEMA_signal_3875, n4190}), .c ({state_out_s1[180], state_out_s0[180]}) ) ;
    xor_HPC2 U4532 ( .a ({new_AGEMA_signal_3477, n4193}), .b ({new_AGEMA_signal_3463, n4192}), .c ({new_AGEMA_signal_3876, n4194}) ) ;
    xnor_HPC2 U4533 ( .a ({new_AGEMA_signal_3460, n4204}), .b ({new_AGEMA_signal_3876, n4194}), .c ({state_out_s1[179], state_out_s0[179]}) ) ;
    xor_HPC2 U4534 ( .a ({new_AGEMA_signal_3458, n4212}), .b ({new_AGEMA_signal_3475, n4195}), .c ({new_AGEMA_signal_3877, n4196}) ) ;
    xnor_HPC2 U4535 ( .a ({new_AGEMA_signal_3460, n4204}), .b ({new_AGEMA_signal_3877, n4196}), .c ({state_out_s1[178], state_out_s0[178]}) ) ;
    xor_HPC2 U4536 ( .a ({new_AGEMA_signal_3458, n4212}), .b ({new_AGEMA_signal_3454, n4213}), .c ({new_AGEMA_signal_3878, n4197}) ) ;
    xnor_HPC2 U4537 ( .a ({new_AGEMA_signal_3472, n4198}), .b ({new_AGEMA_signal_3878, n4197}), .c ({state_out_s1[177], state_out_s0[177]}) ) ;
    xnor_HPC2 U4538 ( .a ({new_AGEMA_signal_3469, n4199}), .b ({new_AGEMA_signal_3454, n4213}), .c ({new_AGEMA_signal_3879, n4200}) ) ;
    xnor_HPC2 U4539 ( .a ({new_AGEMA_signal_3879, n4200}), .b ({new_AGEMA_signal_3507, n4202}), .c ({state_out_s1[176], state_out_s0[176]}) ) ;
    xnor_HPC2 U4540 ( .a ({new_AGEMA_signal_4565, n4219}), .b ({new_AGEMA_signal_3467, n4201}), .c ({new_AGEMA_signal_4607, n4203}) ) ;
    xnor_HPC2 U4541 ( .a ({new_AGEMA_signal_4607, n4203}), .b ({new_AGEMA_signal_3507, n4202}), .c ({state_out_s1[191], state_out_s0[191]}) ) ;
    xnor_HPC2 U4542 ( .a ({new_AGEMA_signal_3460, n4204}), .b ({new_AGEMA_signal_4143, n4228}), .c ({new_AGEMA_signal_4436, n4207}) ) ;
    xnor_HPC2 U4543 ( .a ({1'b0, n4206}), .b ({new_AGEMA_signal_3514, n4205}), .c ({new_AGEMA_signal_3880, n4237}) ) ;
    xnor_HPC2 U4544 ( .a ({new_AGEMA_signal_4436, n4207}), .b ({new_AGEMA_signal_3880, n4237}), .c ({state_out_s1[189], state_out_s0[189]}) ) ;
    xor_HPC2 U4545 ( .a ({new_AGEMA_signal_2843, n4208}), .b ({new_AGEMA_signal_3208, z2[4]}), .c ({new_AGEMA_signal_3516, n4209}) ) ;
    xnor_HPC2 U4546 ( .a ({new_AGEMA_signal_3829, n4210}), .b ({new_AGEMA_signal_3516, n4209}), .c ({new_AGEMA_signal_4195, n4211}) ) ;
    xnor_HPC2 U4547 ( .a ({new_AGEMA_signal_3458, n4212}), .b ({new_AGEMA_signal_4195, n4211}), .c ({state_out_s1[188], state_out_s0[188]}) ) ;
    xnor_HPC2 U4548 ( .a ({new_AGEMA_signal_4564, n4262}), .b ({new_AGEMA_signal_3454, n4213}), .c ({new_AGEMA_signal_4608, n4214}) ) ;
    xnor_HPC2 U4549 ( .a ({new_AGEMA_signal_4608, n4214}), .b ({new_AGEMA_signal_3510, n4250}), .c ({state_out_s1[187], state_out_s0[187]}) ) ;
    xnor_HPC2 U4550 ( .a ({new_AGEMA_signal_3508, n4215}), .b ({new_AGEMA_signal_3505, n4220}), .c ({new_AGEMA_signal_3881, n4216}) ) ;
    xnor_HPC2 U4551 ( .a ({new_AGEMA_signal_3881, n4216}), .b ({new_AGEMA_signal_4138, n4217}), .c ({state_out_s1[132], state_out_s0[132]}) ) ;
    xnor_HPC2 U4552 ( .a ({new_AGEMA_signal_4138, n4217}), .b ({new_AGEMA_signal_3823, n4222}), .c ({new_AGEMA_signal_4439, n4218}) ) ;
    xnor_HPC2 U4553 ( .a ({new_AGEMA_signal_4565, n4219}), .b ({new_AGEMA_signal_4439, n4218}), .c ({state_out_s1[185], state_out_s0[185]}) ) ;
    xor_HPC2 U4554 ( .a ({new_AGEMA_signal_3505, n4220}), .b ({new_AGEMA_signal_3504, n4223}), .c ({new_AGEMA_signal_3882, n4221}) ) ;
    xnor_HPC2 U4555 ( .a ({new_AGEMA_signal_3823, n4222}), .b ({new_AGEMA_signal_3882, n4221}), .c ({state_out_s1[131], state_out_s0[131]}) ) ;
    xor_HPC2 U4556 ( .a ({new_AGEMA_signal_3817, n4224}), .b ({new_AGEMA_signal_3504, n4223}), .c ({new_AGEMA_signal_4197, n4225}) ) ;
    xnor_HPC2 U4557 ( .a ({new_AGEMA_signal_3503, n4226}), .b ({new_AGEMA_signal_4197, n4225}), .c ({state_out_s1[130], state_out_s0[130]}) ) ;
    xor_HPC2 U4558 ( .a ({new_AGEMA_signal_3579, z3[6]}), .b ({state_in_s1[254], state_in_s0[254]}), .c ({new_AGEMA_signal_3883, n4227}) ) ;
    xnor_HPC2 U4559 ( .a ({new_AGEMA_signal_4143, n4228}), .b ({new_AGEMA_signal_3883, n4227}), .c ({new_AGEMA_signal_4441, n4235}) ) ;
    xnor_HPC2 U4560 ( .a ({new_AGEMA_signal_4091, n4230}), .b ({new_AGEMA_signal_4100, n4229}), .c ({new_AGEMA_signal_4442, n4231}) ) ;
    xnor_HPC2 U4561 ( .a ({new_AGEMA_signal_4441, n4235}), .b ({new_AGEMA_signal_4442, n4231}), .c ({state_out_s1[254], state_out_s0[254]}) ) ;
    xnor_HPC2 U4562 ( .a ({new_AGEMA_signal_4123, n4233}), .b ({new_AGEMA_signal_4136, n4232}), .c ({new_AGEMA_signal_4443, n4234}) ) ;
    xnor_HPC2 U4563 ( .a ({new_AGEMA_signal_4441, n4235}), .b ({new_AGEMA_signal_4443, n4234}), .c ({state_out_s1[205], state_out_s0[205]}) ) ;
    xnor_HPC2 U4564 ( .a ({new_AGEMA_signal_4441, n4235}), .b ({new_AGEMA_signal_4092, n4263}), .c ({new_AGEMA_signal_4570, n4236}) ) ;
    xnor_HPC2 U4565 ( .a ({new_AGEMA_signal_4570, n4236}), .b ({new_AGEMA_signal_4130, n4266}), .c ({state_out_s1[196], state_out_s0[196]}) ) ;
    xnor_HPC2 U4566 ( .a ({new_AGEMA_signal_3574, z3[5]}), .b ({state_in_s1[253], state_in_s0[253]}), .c ({new_AGEMA_signal_3884, n4238}) ) ;
    xnor_HPC2 U4567 ( .a ({new_AGEMA_signal_3884, n4238}), .b ({new_AGEMA_signal_3880, n4237}), .c ({new_AGEMA_signal_4198, n4247}) ) ;
    xnor_HPC2 U4568 ( .a ({new_AGEMA_signal_4097, n4239}), .b ({new_AGEMA_signal_4198, n4247}), .c ({new_AGEMA_signal_4444, n4240}) ) ;
    xnor_HPC2 U4569 ( .a ({new_AGEMA_signal_4089, n4241}), .b ({new_AGEMA_signal_4444, n4240}), .c ({state_out_s1[253], state_out_s0[253]}) ) ;
    xnor_HPC2 U4570 ( .a ({new_AGEMA_signal_4122, n4243}), .b ({new_AGEMA_signal_4134, n4242}), .c ({new_AGEMA_signal_4445, n4244}) ) ;
    xnor_HPC2 U4571 ( .a ({new_AGEMA_signal_4445, n4244}), .b ({new_AGEMA_signal_4198, n4247}), .c ({state_out_s1[204], state_out_s0[204]}) ) ;
    xnor_HPC2 U4572 ( .a ({new_AGEMA_signal_4129, n4246}), .b ({new_AGEMA_signal_4088, n4245}), .c ({new_AGEMA_signal_4446, n4248}) ) ;
    xnor_HPC2 U4573 ( .a ({new_AGEMA_signal_4446, n4248}), .b ({new_AGEMA_signal_4198, n4247}), .c ({state_out_s1[195], state_out_s0[195]}) ) ;
    xor_HPC2 U4574 ( .a ({new_AGEMA_signal_3563, z3[4]}), .b ({state_in_s1[252], state_in_s0[252]}), .c ({new_AGEMA_signal_3885, n4249}) ) ;
    xnor_HPC2 U4575 ( .a ({new_AGEMA_signal_3510, n4250}), .b ({new_AGEMA_signal_3885, n4249}), .c ({new_AGEMA_signal_4199, n4260}) ) ;
    xnor_HPC2 U4576 ( .a ({new_AGEMA_signal_4199, n4260}), .b ({new_AGEMA_signal_4121, n4251}), .c ({new_AGEMA_signal_4447, n4252}) ) ;
    xnor_HPC2 U4577 ( .a ({new_AGEMA_signal_4133, n4253}), .b ({new_AGEMA_signal_4447, n4252}), .c ({state_out_s1[203], state_out_s0[203]}) ) ;
    xor_HPC2 U4578 ( .a ({new_AGEMA_signal_4094, n4255}), .b ({new_AGEMA_signal_4086, n4254}), .c ({new_AGEMA_signal_4448, n4256}) ) ;
    xnor_HPC2 U4579 ( .a ({new_AGEMA_signal_4199, n4260}), .b ({new_AGEMA_signal_4448, n4256}), .c ({state_out_s1[252], state_out_s0[252]}) ) ;
    xor_HPC2 U4580 ( .a ({new_AGEMA_signal_4085, n4258}), .b ({new_AGEMA_signal_4128, n4257}), .c ({new_AGEMA_signal_4449, n4259}) ) ;
    xnor_HPC2 U4581 ( .a ({new_AGEMA_signal_4199, n4260}), .b ({new_AGEMA_signal_4449, n4259}), .c ({state_out_s1[194], state_out_s0[194]}) ) ;
    xnor_HPC2 U4582 ( .a ({new_AGEMA_signal_3552, z3[3]}), .b ({state_in_s1[251], state_in_s0[251]}), .c ({new_AGEMA_signal_3886, n4261}) ) ;
    xnor_HPC2 U4583 ( .a ({new_AGEMA_signal_4564, n4262}), .b ({new_AGEMA_signal_3886, n4261}), .c ({new_AGEMA_signal_4611, n4272}) ) ;
    xnor_HPC2 U4584 ( .a ({new_AGEMA_signal_4082, n4264}), .b ({new_AGEMA_signal_4092, n4263}), .c ({new_AGEMA_signal_4450, n4265}) ) ;
    xnor_HPC2 U4585 ( .a ({new_AGEMA_signal_4611, n4272}), .b ({new_AGEMA_signal_4450, n4265}), .c ({state_out_s1[251], state_out_s0[251]}) ) ;
    xnor_HPC2 U4586 ( .a ({new_AGEMA_signal_4120, n4267}), .b ({new_AGEMA_signal_4130, n4266}), .c ({new_AGEMA_signal_4451, n4268}) ) ;
    xnor_HPC2 U4587 ( .a ({new_AGEMA_signal_4611, n4272}), .b ({new_AGEMA_signal_4451, n4268}), .c ({state_out_s1[202], state_out_s0[202]}) ) ;
    xnor_HPC2 U4588 ( .a ({new_AGEMA_signal_4127, n4270}), .b ({new_AGEMA_signal_4083, n4269}), .c ({new_AGEMA_signal_4452, n4271}) ) ;
    xnor_HPC2 U4589 ( .a ({new_AGEMA_signal_4611, n4272}), .b ({new_AGEMA_signal_4452, n4271}), .c ({state_out_s1[193], state_out_s0[193]}) ) ;
    nor_HPC2 SboxInst_U512 ( .a ({new_AGEMA_signal_2989, y2[0]}), .b ({new_AGEMA_signal_2890, SboxInst_n384}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_3517, z1[0]}) ) ;
    nor_HPC2 SboxInst_U511 ( .a ({new_AGEMA_signal_2704, n3290}), .b ({new_AGEMA_signal_2979, SboxInst_n383}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_2991, z1[10]}) ) ;
    nor_HPC2 SboxInst_U510 ( .a ({new_AGEMA_signal_2709, n3289}), .b ({new_AGEMA_signal_2977, SboxInst_n382}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_2992, z1[11]}) ) ;
    nor_HPC2 SboxInst_U509 ( .a ({new_AGEMA_signal_2717, n3288}), .b ({new_AGEMA_signal_2975, SboxInst_n381}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_2993, z1[12]}) ) ;
    nor_HPC2 SboxInst_U508 ( .a ({new_AGEMA_signal_2727, n3286}), .b ({new_AGEMA_signal_2974, SboxInst_n380}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_2994, z1[13]}) ) ;
    nor_HPC2 SboxInst_U507 ( .a ({new_AGEMA_signal_2733, n3285}), .b ({new_AGEMA_signal_2971, SboxInst_n379}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_2995, z1[14]}) ) ;
    nor_HPC2 SboxInst_U506 ( .a ({new_AGEMA_signal_2742, n3284}), .b ({new_AGEMA_signal_2970, SboxInst_n378}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_2996, z1[15]}) ) ;
    nor_HPC2 SboxInst_U505 ( .a ({new_AGEMA_signal_2750, n3283}), .b ({new_AGEMA_signal_2968, SboxInst_n377}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_2997, z1[16]}) ) ;
    nor_HPC2 SboxInst_U504 ( .a ({new_AGEMA_signal_2755, n3282}), .b ({new_AGEMA_signal_2964, SboxInst_n376}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_2998, z1[17]}) ) ;
    nor_HPC2 SboxInst_U503 ( .a ({new_AGEMA_signal_2760, n3281}), .b ({new_AGEMA_signal_2978, SboxInst_n375}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_2999, z1[18]}) ) ;
    nor_HPC2 SboxInst_U502 ( .a ({new_AGEMA_signal_2695, n3280}), .b ({new_AGEMA_signal_2976, SboxInst_n374}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_3000, z1[19]}) ) ;
    nor_HPC2 SboxInst_U501 ( .a ({new_AGEMA_signal_3513, y2[1]}), .b ({new_AGEMA_signal_2896, SboxInst_n373}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_3887, z1[1]}) ) ;
    nor_HPC2 SboxInst_U500 ( .a ({new_AGEMA_signal_2701, n3279}), .b ({new_AGEMA_signal_2973, SboxInst_n372}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_3001, z1[20]}) ) ;
    nor_HPC2 SboxInst_U499 ( .a ({new_AGEMA_signal_2712, n3278}), .b ({new_AGEMA_signal_2972, SboxInst_n371}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_3002, z1[21]}) ) ;
    nor_HPC2 SboxInst_U498 ( .a ({new_AGEMA_signal_2719, n3277}), .b ({new_AGEMA_signal_2969, SboxInst_n370}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_3003, z1[22]}) ) ;
    nor_HPC2 SboxInst_U497 ( .a ({new_AGEMA_signal_2724, n3276}), .b ({new_AGEMA_signal_2967, SboxInst_n369}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_3004, z1[23]}) ) ;
    nor_HPC2 SboxInst_U496 ( .a ({new_AGEMA_signal_2736, n3275}), .b ({new_AGEMA_signal_2965, SboxInst_n368}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_3005, z1[24]}) ) ;
    nor_HPC2 SboxInst_U495 ( .a ({new_AGEMA_signal_2744, n3274}), .b ({new_AGEMA_signal_2980, SboxInst_n367}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_3006, z1[25]}) ) ;
    nor_HPC2 SboxInst_U494 ( .a ({new_AGEMA_signal_2698, n3273}), .b ({new_AGEMA_signal_2987, SboxInst_n366}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_3007, z1[26]}) ) ;
    nor_HPC2 SboxInst_U493 ( .a ({new_AGEMA_signal_2707, n3272}), .b ({new_AGEMA_signal_2985, SboxInst_n365}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_3008, z1[27]}) ) ;
    nor_HPC2 SboxInst_U492 ( .a ({new_AGEMA_signal_2714, n3271}), .b ({new_AGEMA_signal_2984, SboxInst_n364}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_3009, z1[28]}) ) ;
    nor_HPC2 SboxInst_U491 ( .a ({new_AGEMA_signal_2721, n3270}), .b ({new_AGEMA_signal_2983, SboxInst_n363}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_3010, z1[29]}) ) ;
    nor_HPC2 SboxInst_U490 ( .a ({new_AGEMA_signal_3824, n3287}), .b ({new_AGEMA_signal_2895, SboxInst_n362}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_4200, z1[2]}) ) ;
    nor_HPC2 SboxInst_U489 ( .a ({new_AGEMA_signal_2730, n3269}), .b ({new_AGEMA_signal_2982, SboxInst_n361}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_3011, z1[30]}) ) ;
    nor_HPC2 SboxInst_U488 ( .a ({new_AGEMA_signal_2739, n3268}), .b ({new_AGEMA_signal_2981, SboxInst_n360}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_3012, z1[31]}) ) ;
    nor_HPC2 SboxInst_U487 ( .a ({new_AGEMA_signal_2747, n3267}), .b ({new_AGEMA_signal_2872, SboxInst_n359}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_3013, z1[32]}) ) ;
    nor_HPC2 SboxInst_U486 ( .a ({new_AGEMA_signal_2753, n3266}), .b ({new_AGEMA_signal_2871, SboxInst_n358}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_3014, z1[33]}) ) ;
    nor_HPC2 SboxInst_U485 ( .a ({new_AGEMA_signal_2758, n3265}), .b ({new_AGEMA_signal_2870, SboxInst_n357}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_3015, z1[34]}) ) ;
    nor_HPC2 SboxInst_U484 ( .a ({new_AGEMA_signal_2763, n3264}), .b ({new_AGEMA_signal_2869, SboxInst_n356}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_3016, z1[35]}) ) ;
    nor_HPC2 SboxInst_U483 ( .a ({new_AGEMA_signal_2766, n3263}), .b ({new_AGEMA_signal_2867, SboxInst_n355}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_3017, z1[36]}) ) ;
    nor_HPC2 SboxInst_U482 ( .a ({new_AGEMA_signal_2769, n3262}), .b ({new_AGEMA_signal_2865, SboxInst_n354}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_3018, z1[37]}) ) ;
    nor_HPC2 SboxInst_U481 ( .a ({new_AGEMA_signal_2772, n3261}), .b ({new_AGEMA_signal_2863, SboxInst_n353}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_3019, z1[38]}) ) ;
    nor_HPC2 SboxInst_U480 ( .a ({new_AGEMA_signal_2775, n3260}), .b ({new_AGEMA_signal_2860, SboxInst_n352}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_3020, z1[39]}) ) ;
    nor_HPC2 SboxInst_U479 ( .a ({new_AGEMA_signal_4432, n3233}), .b ({new_AGEMA_signal_2894, SboxInst_n351}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_4577, z1[3]}) ) ;
    nor_HPC2 SboxInst_U478 ( .a ({new_AGEMA_signal_2778, n3259}), .b ({new_AGEMA_signal_2861, SboxInst_n350}), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_3021, z1[40]}) ) ;
    nor_HPC2 SboxInst_U477 ( .a ({new_AGEMA_signal_2780, n3258}), .b ({new_AGEMA_signal_2868, SboxInst_n349}), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_3022, z1[41]}) ) ;
    nor_HPC2 SboxInst_U476 ( .a ({new_AGEMA_signal_2783, n3257}), .b ({new_AGEMA_signal_2866, SboxInst_n348}), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_3023, z1[42]}) ) ;
    nor_HPC2 SboxInst_U475 ( .a ({new_AGEMA_signal_2786, n3256}), .b ({new_AGEMA_signal_2864, SboxInst_n347}), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_3024, z1[43]}) ) ;
    nor_HPC2 SboxInst_U474 ( .a ({new_AGEMA_signal_2788, n3255}), .b ({new_AGEMA_signal_2862, SboxInst_n346}), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_3025, z1[44]}) ) ;
    nor_HPC2 SboxInst_U473 ( .a ({new_AGEMA_signal_2790, n3254}), .b ({new_AGEMA_signal_2859, SboxInst_n345}), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_3026, z1[45]}) ) ;
    nor_HPC2 SboxInst_U472 ( .a ({new_AGEMA_signal_2793, n3253}), .b ({new_AGEMA_signal_2877, SboxInst_n344}), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_3027, z1[46]}) ) ;
    nor_HPC2 SboxInst_U471 ( .a ({new_AGEMA_signal_2795, n3252}), .b ({new_AGEMA_signal_2875, SboxInst_n343}), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_3028, z1[47]}) ) ;
    nor_HPC2 SboxInst_U470 ( .a ({new_AGEMA_signal_2797, n3251}), .b ({new_AGEMA_signal_2873, SboxInst_n342}), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_3029, z1[48]}) ) ;
    nor_HPC2 SboxInst_U469 ( .a ({new_AGEMA_signal_2800, n3250}), .b ({new_AGEMA_signal_2880, SboxInst_n341}), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_3030, z1[49]}) ) ;
    nor_HPC2 SboxInst_U468 ( .a ({new_AGEMA_signal_2990, n3232}), .b ({new_AGEMA_signal_2892, SboxInst_n340}), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_3518, z1[4]}) ) ;
    nor_HPC2 SboxInst_U467 ( .a ({new_AGEMA_signal_2803, n3249}), .b ({new_AGEMA_signal_2879, SboxInst_n339}), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_3031, z1[50]}) ) ;
    nor_HPC2 SboxInst_U466 ( .a ({new_AGEMA_signal_2805, n3248}), .b ({new_AGEMA_signal_2878, SboxInst_n338}), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_3032, z1[51]}) ) ;
    nor_HPC2 SboxInst_U465 ( .a ({new_AGEMA_signal_2807, n3247}), .b ({new_AGEMA_signal_2876, SboxInst_n337}), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_3033, z1[52]}) ) ;
    nor_HPC2 SboxInst_U464 ( .a ({new_AGEMA_signal_2810, n3246}), .b ({new_AGEMA_signal_2874, SboxInst_n336}), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_3034, z1[53]}) ) ;
    nor_HPC2 SboxInst_U463 ( .a ({new_AGEMA_signal_2813, n3245}), .b ({new_AGEMA_signal_2884, SboxInst_n335}), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_3035, z1[54]}) ) ;
    nor_HPC2 SboxInst_U462 ( .a ({new_AGEMA_signal_2816, n3244}), .b ({new_AGEMA_signal_2881, SboxInst_n334}), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_3036, z1[55]}) ) ;
    nor_HPC2 SboxInst_U461 ( .a ({new_AGEMA_signal_2819, n3243}), .b ({new_AGEMA_signal_2883, SboxInst_n333}), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_3037, z1[56]}) ) ;
    nor_HPC2 SboxInst_U460 ( .a ({new_AGEMA_signal_2821, n3242}), .b ({new_AGEMA_signal_2888, SboxInst_n332}), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_3038, z1[57]}) ) ;
    nor_HPC2 SboxInst_U459 ( .a ({new_AGEMA_signal_2823, n3241}), .b ({new_AGEMA_signal_2887, SboxInst_n331}), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_3039, z1[58]}) ) ;
    nor_HPC2 SboxInst_U458 ( .a ({new_AGEMA_signal_2825, n3240}), .b ({new_AGEMA_signal_2886, SboxInst_n330}), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_3040, z1[59]}) ) ;
    nor_HPC2 SboxInst_U457 ( .a ({new_AGEMA_signal_3515, n3231}), .b ({new_AGEMA_signal_2891, SboxInst_n329}), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_3888, z1[5]}) ) ;
    nor_HPC2 SboxInst_U456 ( .a ({new_AGEMA_signal_2828, n3238}), .b ({new_AGEMA_signal_2885, SboxInst_n328}), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_3041, z1[60]}) ) ;
    nor_HPC2 SboxInst_U455 ( .a ({new_AGEMA_signal_2837, n3236}), .b ({new_AGEMA_signal_2882, SboxInst_n327}), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_3042, z1[61]}) ) ;
    nor_HPC2 SboxInst_U454 ( .a ({new_AGEMA_signal_2840, n3235}), .b ({new_AGEMA_signal_2893, SboxInst_n326}), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_3043, z1[62]}) ) ;
    nor_HPC2 SboxInst_U453 ( .a ({new_AGEMA_signal_2846, n3234}), .b ({new_AGEMA_signal_2889, SboxInst_n325}), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_3044, z1[63]}) ) ;
    nor_HPC2 SboxInst_U452 ( .a ({new_AGEMA_signal_3826, n3230}), .b ({new_AGEMA_signal_2966, SboxInst_n324}), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_4201, z1[6]}) ) ;
    nor_HPC2 SboxInst_U451 ( .a ({new_AGEMA_signal_4433, n3239}), .b ({new_AGEMA_signal_2963, SboxInst_n323}), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_4578, z1[7]}) ) ;
    nor_HPC2 SboxInst_U450 ( .a ({new_AGEMA_signal_2834, n3237}), .b ({new_AGEMA_signal_2988, SboxInst_n322}), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_3045, z1[8]}) ) ;
    nor_HPC2 SboxInst_U449 ( .a ({new_AGEMA_signal_2692, n3291}), .b ({new_AGEMA_signal_2986, SboxInst_n321}), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_3046, z1[9]}) ) ;
    nor_HPC2 SboxInst_U448 ( .a ({new_AGEMA_signal_2527, y4[0]}), .b ({new_AGEMA_signal_3047, SboxInst_n320}), .clk (clk), .r (Fresh[64]), .c ({new_AGEMA_signal_3519, z3[0]}) ) ;
    nor_HPC2 SboxInst_U446 ( .a ({new_AGEMA_signal_2524, y4[10]}), .b ({new_AGEMA_signal_3048, SboxInst_n319}), .clk (clk), .r (Fresh[65]), .c ({new_AGEMA_signal_3520, z3[10]}) ) ;
    nor_HPC2 SboxInst_U444 ( .a ({new_AGEMA_signal_2521, y4[11]}), .b ({new_AGEMA_signal_3049, SboxInst_n318}), .clk (clk), .r (Fresh[66]), .c ({new_AGEMA_signal_3521, z3[11]}) ) ;
    nor_HPC2 SboxInst_U442 ( .a ({new_AGEMA_signal_2518, y4[12]}), .b ({new_AGEMA_signal_3050, SboxInst_n317}), .clk (clk), .r (Fresh[67]), .c ({new_AGEMA_signal_3522, z3[12]}) ) ;
    nor_HPC2 SboxInst_U440 ( .a ({new_AGEMA_signal_2515, y4[13]}), .b ({new_AGEMA_signal_3051, SboxInst_n316}), .clk (clk), .r (Fresh[68]), .c ({new_AGEMA_signal_3523, z3[13]}) ) ;
    nor_HPC2 SboxInst_U438 ( .a ({new_AGEMA_signal_2512, y4[14]}), .b ({new_AGEMA_signal_3052, SboxInst_n315}), .clk (clk), .r (Fresh[69]), .c ({new_AGEMA_signal_3524, z3[14]}) ) ;
    nor_HPC2 SboxInst_U436 ( .a ({new_AGEMA_signal_2509, y4[15]}), .b ({new_AGEMA_signal_3053, SboxInst_n314}), .clk (clk), .r (Fresh[70]), .c ({new_AGEMA_signal_3525, z3[15]}) ) ;
    nor_HPC2 SboxInst_U434 ( .a ({new_AGEMA_signal_2506, y4[16]}), .b ({new_AGEMA_signal_3054, SboxInst_n313}), .clk (clk), .r (Fresh[71]), .c ({new_AGEMA_signal_3526, z3[16]}) ) ;
    nor_HPC2 SboxInst_U432 ( .a ({new_AGEMA_signal_2503, y4[17]}), .b ({new_AGEMA_signal_3055, SboxInst_n312}), .clk (clk), .r (Fresh[72]), .c ({new_AGEMA_signal_3527, z3[17]}) ) ;
    nor_HPC2 SboxInst_U430 ( .a ({new_AGEMA_signal_2500, y4[18]}), .b ({new_AGEMA_signal_3056, SboxInst_n311}), .clk (clk), .r (Fresh[73]), .c ({new_AGEMA_signal_3528, z3[18]}) ) ;
    nor_HPC2 SboxInst_U428 ( .a ({new_AGEMA_signal_2497, y4[19]}), .b ({new_AGEMA_signal_3057, SboxInst_n310}), .clk (clk), .r (Fresh[74]), .c ({new_AGEMA_signal_3529, z3[19]}) ) ;
    nor_HPC2 SboxInst_U426 ( .a ({new_AGEMA_signal_2494, y4[1]}), .b ({new_AGEMA_signal_3058, SboxInst_n309}), .clk (clk), .r (Fresh[75]), .c ({new_AGEMA_signal_3530, z3[1]}) ) ;
    nor_HPC2 SboxInst_U424 ( .a ({new_AGEMA_signal_2491, y4[20]}), .b ({new_AGEMA_signal_3059, SboxInst_n308}), .clk (clk), .r (Fresh[76]), .c ({new_AGEMA_signal_3531, z3[20]}) ) ;
    nor_HPC2 SboxInst_U422 ( .a ({new_AGEMA_signal_2488, y4[21]}), .b ({new_AGEMA_signal_3060, SboxInst_n307}), .clk (clk), .r (Fresh[77]), .c ({new_AGEMA_signal_3532, z3[21]}) ) ;
    nor_HPC2 SboxInst_U420 ( .a ({new_AGEMA_signal_2485, y4[22]}), .b ({new_AGEMA_signal_3061, SboxInst_n306}), .clk (clk), .r (Fresh[78]), .c ({new_AGEMA_signal_3533, z3[22]}) ) ;
    nor_HPC2 SboxInst_U418 ( .a ({new_AGEMA_signal_2482, y4[23]}), .b ({new_AGEMA_signal_3062, SboxInst_n305}), .clk (clk), .r (Fresh[79]), .c ({new_AGEMA_signal_3534, z3[23]}) ) ;
    nor_HPC2 SboxInst_U416 ( .a ({new_AGEMA_signal_2479, y4[24]}), .b ({new_AGEMA_signal_3063, SboxInst_n304}), .clk (clk), .r (Fresh[80]), .c ({new_AGEMA_signal_3535, z3[24]}) ) ;
    nor_HPC2 SboxInst_U414 ( .a ({new_AGEMA_signal_2476, y4[25]}), .b ({new_AGEMA_signal_3064, SboxInst_n303}), .clk (clk), .r (Fresh[81]), .c ({new_AGEMA_signal_3536, z3[25]}) ) ;
    nor_HPC2 SboxInst_U412 ( .a ({new_AGEMA_signal_2473, y4[26]}), .b ({new_AGEMA_signal_3065, SboxInst_n302}), .clk (clk), .r (Fresh[82]), .c ({new_AGEMA_signal_3537, z3[26]}) ) ;
    nor_HPC2 SboxInst_U410 ( .a ({new_AGEMA_signal_2470, y4[27]}), .b ({new_AGEMA_signal_3066, SboxInst_n301}), .clk (clk), .r (Fresh[83]), .c ({new_AGEMA_signal_3538, z3[27]}) ) ;
    nor_HPC2 SboxInst_U408 ( .a ({new_AGEMA_signal_2467, y4[28]}), .b ({new_AGEMA_signal_3067, SboxInst_n300}), .clk (clk), .r (Fresh[84]), .c ({new_AGEMA_signal_3539, z3[28]}) ) ;
    nor_HPC2 SboxInst_U406 ( .a ({new_AGEMA_signal_2464, y4[29]}), .b ({new_AGEMA_signal_3068, SboxInst_n299}), .clk (clk), .r (Fresh[85]), .c ({new_AGEMA_signal_3540, z3[29]}) ) ;
    nor_HPC2 SboxInst_U404 ( .a ({new_AGEMA_signal_2461, y4[2]}), .b ({new_AGEMA_signal_3069, SboxInst_n298}), .clk (clk), .r (Fresh[86]), .c ({new_AGEMA_signal_3541, z3[2]}) ) ;
    nor_HPC2 SboxInst_U402 ( .a ({new_AGEMA_signal_2458, y4[30]}), .b ({new_AGEMA_signal_3070, SboxInst_n297}), .clk (clk), .r (Fresh[87]), .c ({new_AGEMA_signal_3542, z3[30]}) ) ;
    nor_HPC2 SboxInst_U400 ( .a ({new_AGEMA_signal_2455, y4[31]}), .b ({new_AGEMA_signal_3071, SboxInst_n296}), .clk (clk), .r (Fresh[88]), .c ({new_AGEMA_signal_3543, z3[31]}) ) ;
    nor_HPC2 SboxInst_U398 ( .a ({new_AGEMA_signal_2452, y4[32]}), .b ({new_AGEMA_signal_3072, SboxInst_n295}), .clk (clk), .r (Fresh[89]), .c ({new_AGEMA_signal_3544, z3[32]}) ) ;
    nor_HPC2 SboxInst_U396 ( .a ({new_AGEMA_signal_2449, y4[33]}), .b ({new_AGEMA_signal_3073, SboxInst_n294}), .clk (clk), .r (Fresh[90]), .c ({new_AGEMA_signal_3545, z3[33]}) ) ;
    nor_HPC2 SboxInst_U394 ( .a ({new_AGEMA_signal_2446, y4[34]}), .b ({new_AGEMA_signal_3074, SboxInst_n293}), .clk (clk), .r (Fresh[91]), .c ({new_AGEMA_signal_3546, z3[34]}) ) ;
    nor_HPC2 SboxInst_U392 ( .a ({new_AGEMA_signal_2443, y4[35]}), .b ({new_AGEMA_signal_3075, SboxInst_n292}), .clk (clk), .r (Fresh[92]), .c ({new_AGEMA_signal_3547, z3[35]}) ) ;
    nor_HPC2 SboxInst_U390 ( .a ({new_AGEMA_signal_2440, y4[36]}), .b ({new_AGEMA_signal_3076, SboxInst_n291}), .clk (clk), .r (Fresh[93]), .c ({new_AGEMA_signal_3548, z3[36]}) ) ;
    nor_HPC2 SboxInst_U388 ( .a ({new_AGEMA_signal_2437, y4[37]}), .b ({new_AGEMA_signal_3077, SboxInst_n290}), .clk (clk), .r (Fresh[94]), .c ({new_AGEMA_signal_3549, z3[37]}) ) ;
    nor_HPC2 SboxInst_U386 ( .a ({new_AGEMA_signal_2434, y4[38]}), .b ({new_AGEMA_signal_3078, SboxInst_n289}), .clk (clk), .r (Fresh[95]), .c ({new_AGEMA_signal_3550, z3[38]}) ) ;
    nor_HPC2 SboxInst_U384 ( .a ({new_AGEMA_signal_2431, y4[39]}), .b ({new_AGEMA_signal_3079, SboxInst_n288}), .clk (clk), .r (Fresh[96]), .c ({new_AGEMA_signal_3551, z3[39]}) ) ;
    nor_HPC2 SboxInst_U382 ( .a ({new_AGEMA_signal_2428, y4[3]}), .b ({new_AGEMA_signal_3080, SboxInst_n287}), .clk (clk), .r (Fresh[97]), .c ({new_AGEMA_signal_3552, z3[3]}) ) ;
    nor_HPC2 SboxInst_U380 ( .a ({new_AGEMA_signal_2425, y4[40]}), .b ({new_AGEMA_signal_3081, SboxInst_n286}), .clk (clk), .r (Fresh[98]), .c ({new_AGEMA_signal_3553, z3[40]}) ) ;
    nor_HPC2 SboxInst_U378 ( .a ({new_AGEMA_signal_2422, y4[41]}), .b ({new_AGEMA_signal_3082, SboxInst_n285}), .clk (clk), .r (Fresh[99]), .c ({new_AGEMA_signal_3554, z3[41]}) ) ;
    nor_HPC2 SboxInst_U376 ( .a ({new_AGEMA_signal_2419, y4[42]}), .b ({new_AGEMA_signal_3083, SboxInst_n284}), .clk (clk), .r (Fresh[100]), .c ({new_AGEMA_signal_3555, z3[42]}) ) ;
    nor_HPC2 SboxInst_U374 ( .a ({new_AGEMA_signal_2416, y4[43]}), .b ({new_AGEMA_signal_3084, SboxInst_n283}), .clk (clk), .r (Fresh[101]), .c ({new_AGEMA_signal_3556, z3[43]}) ) ;
    nor_HPC2 SboxInst_U372 ( .a ({new_AGEMA_signal_2413, y4[44]}), .b ({new_AGEMA_signal_3085, SboxInst_n282}), .clk (clk), .r (Fresh[102]), .c ({new_AGEMA_signal_3557, z3[44]}) ) ;
    nor_HPC2 SboxInst_U370 ( .a ({new_AGEMA_signal_2410, y4[45]}), .b ({new_AGEMA_signal_3086, SboxInst_n281}), .clk (clk), .r (Fresh[103]), .c ({new_AGEMA_signal_3558, z3[45]}) ) ;
    nor_HPC2 SboxInst_U368 ( .a ({new_AGEMA_signal_2407, y4[46]}), .b ({new_AGEMA_signal_3087, SboxInst_n280}), .clk (clk), .r (Fresh[104]), .c ({new_AGEMA_signal_3559, z3[46]}) ) ;
    nor_HPC2 SboxInst_U366 ( .a ({new_AGEMA_signal_2404, y4[47]}), .b ({new_AGEMA_signal_3088, SboxInst_n279}), .clk (clk), .r (Fresh[105]), .c ({new_AGEMA_signal_3560, z3[47]}) ) ;
    nor_HPC2 SboxInst_U364 ( .a ({new_AGEMA_signal_2401, y4[48]}), .b ({new_AGEMA_signal_3089, SboxInst_n278}), .clk (clk), .r (Fresh[106]), .c ({new_AGEMA_signal_3561, z3[48]}) ) ;
    nor_HPC2 SboxInst_U362 ( .a ({new_AGEMA_signal_2398, y4[49]}), .b ({new_AGEMA_signal_3090, SboxInst_n277}), .clk (clk), .r (Fresh[107]), .c ({new_AGEMA_signal_3562, z3[49]}) ) ;
    nor_HPC2 SboxInst_U360 ( .a ({new_AGEMA_signal_2395, y4[4]}), .b ({new_AGEMA_signal_3091, SboxInst_n276}), .clk (clk), .r (Fresh[108]), .c ({new_AGEMA_signal_3563, z3[4]}) ) ;
    nor_HPC2 SboxInst_U358 ( .a ({new_AGEMA_signal_2392, y4[50]}), .b ({new_AGEMA_signal_3092, SboxInst_n275}), .clk (clk), .r (Fresh[109]), .c ({new_AGEMA_signal_3564, z3[50]}) ) ;
    nor_HPC2 SboxInst_U356 ( .a ({new_AGEMA_signal_2389, y4[51]}), .b ({new_AGEMA_signal_3093, SboxInst_n274}), .clk (clk), .r (Fresh[110]), .c ({new_AGEMA_signal_3565, z3[51]}) ) ;
    nor_HPC2 SboxInst_U354 ( .a ({new_AGEMA_signal_2386, y4[52]}), .b ({new_AGEMA_signal_3094, SboxInst_n273}), .clk (clk), .r (Fresh[111]), .c ({new_AGEMA_signal_3566, z3[52]}) ) ;
    nor_HPC2 SboxInst_U352 ( .a ({new_AGEMA_signal_2383, y4[53]}), .b ({new_AGEMA_signal_3095, SboxInst_n272}), .clk (clk), .r (Fresh[112]), .c ({new_AGEMA_signal_3567, z3[53]}) ) ;
    nor_HPC2 SboxInst_U350 ( .a ({new_AGEMA_signal_2380, y4[54]}), .b ({new_AGEMA_signal_3096, SboxInst_n271}), .clk (clk), .r (Fresh[113]), .c ({new_AGEMA_signal_3568, z3[54]}) ) ;
    nor_HPC2 SboxInst_U348 ( .a ({new_AGEMA_signal_2377, y4[55]}), .b ({new_AGEMA_signal_3097, SboxInst_n270}), .clk (clk), .r (Fresh[114]), .c ({new_AGEMA_signal_3569, z3[55]}) ) ;
    nor_HPC2 SboxInst_U346 ( .a ({new_AGEMA_signal_2374, y4[56]}), .b ({new_AGEMA_signal_3098, SboxInst_n269}), .clk (clk), .r (Fresh[115]), .c ({new_AGEMA_signal_3570, z3[56]}) ) ;
    nor_HPC2 SboxInst_U344 ( .a ({new_AGEMA_signal_2371, y4[57]}), .b ({new_AGEMA_signal_3099, SboxInst_n268}), .clk (clk), .r (Fresh[116]), .c ({new_AGEMA_signal_3571, z3[57]}) ) ;
    nor_HPC2 SboxInst_U342 ( .a ({new_AGEMA_signal_2368, y4[58]}), .b ({new_AGEMA_signal_3100, SboxInst_n267}), .clk (clk), .r (Fresh[117]), .c ({new_AGEMA_signal_3572, z3[58]}) ) ;
    nor_HPC2 SboxInst_U340 ( .a ({new_AGEMA_signal_2365, y4[59]}), .b ({new_AGEMA_signal_3101, SboxInst_n266}), .clk (clk), .r (Fresh[118]), .c ({new_AGEMA_signal_3573, z3[59]}) ) ;
    nor_HPC2 SboxInst_U338 ( .a ({new_AGEMA_signal_2362, y4[5]}), .b ({new_AGEMA_signal_3102, SboxInst_n265}), .clk (clk), .r (Fresh[119]), .c ({new_AGEMA_signal_3574, z3[5]}) ) ;
    nor_HPC2 SboxInst_U336 ( .a ({new_AGEMA_signal_2359, y4[60]}), .b ({new_AGEMA_signal_3103, SboxInst_n264}), .clk (clk), .r (Fresh[120]), .c ({new_AGEMA_signal_3575, z3[60]}) ) ;
    nor_HPC2 SboxInst_U334 ( .a ({new_AGEMA_signal_2356, y4[61]}), .b ({new_AGEMA_signal_3104, SboxInst_n263}), .clk (clk), .r (Fresh[121]), .c ({new_AGEMA_signal_3576, z3[61]}) ) ;
    nor_HPC2 SboxInst_U332 ( .a ({new_AGEMA_signal_2353, y4[62]}), .b ({new_AGEMA_signal_3105, SboxInst_n262}), .clk (clk), .r (Fresh[122]), .c ({new_AGEMA_signal_3577, z3[62]}) ) ;
    nor_HPC2 SboxInst_U330 ( .a ({new_AGEMA_signal_2350, y4[63]}), .b ({new_AGEMA_signal_3106, SboxInst_n261}), .clk (clk), .r (Fresh[123]), .c ({new_AGEMA_signal_3578, z3[63]}) ) ;
    nor_HPC2 SboxInst_U328 ( .a ({new_AGEMA_signal_2347, y4[6]}), .b ({new_AGEMA_signal_3107, SboxInst_n260}), .clk (clk), .r (Fresh[124]), .c ({new_AGEMA_signal_3579, z3[6]}) ) ;
    nor_HPC2 SboxInst_U326 ( .a ({new_AGEMA_signal_2344, y4[7]}), .b ({new_AGEMA_signal_3108, SboxInst_n259}), .clk (clk), .r (Fresh[125]), .c ({new_AGEMA_signal_3580, z3[7]}) ) ;
    nor_HPC2 SboxInst_U324 ( .a ({new_AGEMA_signal_2341, y4[8]}), .b ({new_AGEMA_signal_3109, SboxInst_n258}), .clk (clk), .r (Fresh[126]), .c ({new_AGEMA_signal_3581, z3[8]}) ) ;
    nor_HPC2 SboxInst_U322 ( .a ({new_AGEMA_signal_2338, y4[9]}), .b ({new_AGEMA_signal_3110, SboxInst_n257}), .clk (clk), .r (Fresh[127]), .c ({new_AGEMA_signal_3582, z3[9]}) ) ;
    nor_HPC2 SboxInst_U320 ( .a ({new_AGEMA_signal_2655, y0[0]}), .b ({new_AGEMA_signal_2911, SboxInst_n256}), .clk (clk), .r (Fresh[128]), .c ({new_AGEMA_signal_3111, z4[0]}) ) ;
    nor_HPC2 SboxInst_U319 ( .a ({new_AGEMA_signal_2653, y0[10]}), .b ({new_AGEMA_signal_2924, SboxInst_n255}), .clk (clk), .r (Fresh[129]), .c ({new_AGEMA_signal_3112, z4[10]}) ) ;
    nor_HPC2 SboxInst_U318 ( .a ({new_AGEMA_signal_2651, y0[11]}), .b ({new_AGEMA_signal_2921, SboxInst_n254}), .clk (clk), .r (Fresh[130]), .c ({new_AGEMA_signal_3113, z4[11]}) ) ;
    nor_HPC2 SboxInst_U317 ( .a ({new_AGEMA_signal_2649, y0[12]}), .b ({new_AGEMA_signal_2919, SboxInst_n253}), .clk (clk), .r (Fresh[131]), .c ({new_AGEMA_signal_3114, z4[12]}) ) ;
    nor_HPC2 SboxInst_U316 ( .a ({new_AGEMA_signal_2647, y0[13]}), .b ({new_AGEMA_signal_2925, SboxInst_n252}), .clk (clk), .r (Fresh[132]), .c ({new_AGEMA_signal_3115, z4[13]}) ) ;
    nor_HPC2 SboxInst_U315 ( .a ({new_AGEMA_signal_2645, y0[14]}), .b ({new_AGEMA_signal_2922, SboxInst_n251}), .clk (clk), .r (Fresh[133]), .c ({new_AGEMA_signal_3116, z4[14]}) ) ;
    nor_HPC2 SboxInst_U314 ( .a ({new_AGEMA_signal_2643, y0[15]}), .b ({new_AGEMA_signal_2918, SboxInst_n250}), .clk (clk), .r (Fresh[134]), .c ({new_AGEMA_signal_3117, z4[15]}) ) ;
    nor_HPC2 SboxInst_U313 ( .a ({new_AGEMA_signal_2641, y0[16]}), .b ({new_AGEMA_signal_2944, SboxInst_n249}), .clk (clk), .r (Fresh[135]), .c ({new_AGEMA_signal_3118, z4[16]}) ) ;
    nor_HPC2 SboxInst_U312 ( .a ({new_AGEMA_signal_2639, y0[17]}), .b ({new_AGEMA_signal_2942, SboxInst_n248}), .clk (clk), .r (Fresh[136]), .c ({new_AGEMA_signal_3119, z4[17]}) ) ;
    nor_HPC2 SboxInst_U311 ( .a ({new_AGEMA_signal_2637, y0[18]}), .b ({new_AGEMA_signal_2940, SboxInst_n247}), .clk (clk), .r (Fresh[137]), .c ({new_AGEMA_signal_3120, z4[18]}) ) ;
    nor_HPC2 SboxInst_U310 ( .a ({new_AGEMA_signal_2635, y0[19]}), .b ({new_AGEMA_signal_2936, SboxInst_n246}), .clk (clk), .r (Fresh[138]), .c ({new_AGEMA_signal_3121, z4[19]}) ) ;
    nor_HPC2 SboxInst_U309 ( .a ({new_AGEMA_signal_2633, y0[1]}), .b ({new_AGEMA_signal_2909, SboxInst_n245}), .clk (clk), .r (Fresh[139]), .c ({new_AGEMA_signal_3122, z4[1]}) ) ;
    nor_HPC2 SboxInst_U308 ( .a ({new_AGEMA_signal_2631, y0[20]}), .b ({new_AGEMA_signal_2934, SboxInst_n244}), .clk (clk), .r (Fresh[140]), .c ({new_AGEMA_signal_3123, z4[20]}) ) ;
    nor_HPC2 SboxInst_U307 ( .a ({new_AGEMA_signal_2629, y0[21]}), .b ({new_AGEMA_signal_2939, SboxInst_n243}), .clk (clk), .r (Fresh[141]), .c ({new_AGEMA_signal_3124, z4[21]}) ) ;
    nor_HPC2 SboxInst_U306 ( .a ({new_AGEMA_signal_2627, y0[22]}), .b ({new_AGEMA_signal_2937, SboxInst_n242}), .clk (clk), .r (Fresh[142]), .c ({new_AGEMA_signal_3125, z4[22]}) ) ;
    nor_HPC2 SboxInst_U305 ( .a ({new_AGEMA_signal_2625, y0[23]}), .b ({new_AGEMA_signal_2935, SboxInst_n241}), .clk (clk), .r (Fresh[143]), .c ({new_AGEMA_signal_3126, z4[23]}) ) ;
    nor_HPC2 SboxInst_U304 ( .a ({new_AGEMA_signal_2623, y0[24]}), .b ({new_AGEMA_signal_2955, SboxInst_n240}), .clk (clk), .r (Fresh[144]), .c ({new_AGEMA_signal_3127, z4[24]}) ) ;
    nor_HPC2 SboxInst_U303 ( .a ({new_AGEMA_signal_2621, y0[25]}), .b ({new_AGEMA_signal_2954, SboxInst_n239}), .clk (clk), .r (Fresh[145]), .c ({new_AGEMA_signal_3128, z4[25]}) ) ;
    nor_HPC2 SboxInst_U302 ( .a ({new_AGEMA_signal_2619, y0[26]}), .b ({new_AGEMA_signal_2952, SboxInst_n238}), .clk (clk), .r (Fresh[146]), .c ({new_AGEMA_signal_3129, z4[26]}) ) ;
    nor_HPC2 SboxInst_U301 ( .a ({new_AGEMA_signal_2617, y0[27]}), .b ({new_AGEMA_signal_2951, SboxInst_n237}), .clk (clk), .r (Fresh[147]), .c ({new_AGEMA_signal_3130, z4[27]}) ) ;
    nor_HPC2 SboxInst_U300 ( .a ({new_AGEMA_signal_2615, y0[28]}), .b ({new_AGEMA_signal_2949, SboxInst_n236}), .clk (clk), .r (Fresh[148]), .c ({new_AGEMA_signal_3131, z4[28]}) ) ;
    nor_HPC2 SboxInst_U299 ( .a ({new_AGEMA_signal_2613, y0[29]}), .b ({new_AGEMA_signal_2953, SboxInst_n235}), .clk (clk), .r (Fresh[149]), .c ({new_AGEMA_signal_3132, z4[29]}) ) ;
    nor_HPC2 SboxInst_U298 ( .a ({new_AGEMA_signal_2611, y0[2]}), .b ({new_AGEMA_signal_2906, SboxInst_n234}), .clk (clk), .r (Fresh[150]), .c ({new_AGEMA_signal_3133, z4[2]}) ) ;
    nor_HPC2 SboxInst_U297 ( .a ({new_AGEMA_signal_2609, y0[30]}), .b ({new_AGEMA_signal_2950, SboxInst_n233}), .clk (clk), .r (Fresh[151]), .c ({new_AGEMA_signal_3134, z4[30]}) ) ;
    nor_HPC2 SboxInst_U296 ( .a ({new_AGEMA_signal_2607, y0[31]}), .b ({new_AGEMA_signal_2948, SboxInst_n232}), .clk (clk), .r (Fresh[152]), .c ({new_AGEMA_signal_3135, z4[31]}) ) ;
    nor_HPC2 SboxInst_U295 ( .a ({new_AGEMA_signal_2605, y0[32]}), .b ({new_AGEMA_signal_2962, SboxInst_n231}), .clk (clk), .r (Fresh[153]), .c ({new_AGEMA_signal_3136, z4[32]}) ) ;
    nor_HPC2 SboxInst_U294 ( .a ({new_AGEMA_signal_2603, y0[33]}), .b ({new_AGEMA_signal_2961, SboxInst_n230}), .clk (clk), .r (Fresh[154]), .c ({new_AGEMA_signal_3137, z4[33]}) ) ;
    nor_HPC2 SboxInst_U293 ( .a ({new_AGEMA_signal_2601, y0[34]}), .b ({new_AGEMA_signal_2959, SboxInst_n229}), .clk (clk), .r (Fresh[155]), .c ({new_AGEMA_signal_3138, z4[34]}) ) ;
    nor_HPC2 SboxInst_U292 ( .a ({new_AGEMA_signal_2599, y0[35]}), .b ({new_AGEMA_signal_2957, SboxInst_n228}), .clk (clk), .r (Fresh[156]), .c ({new_AGEMA_signal_3139, z4[35]}) ) ;
    nor_HPC2 SboxInst_U291 ( .a ({new_AGEMA_signal_2597, y0[36]}), .b ({new_AGEMA_signal_2956, SboxInst_n227}), .clk (clk), .r (Fresh[157]), .c ({new_AGEMA_signal_3140, z4[36]}) ) ;
    nor_HPC2 SboxInst_U290 ( .a ({new_AGEMA_signal_2595, y0[37]}), .b ({new_AGEMA_signal_2960, SboxInst_n226}), .clk (clk), .r (Fresh[158]), .c ({new_AGEMA_signal_3141, z4[37]}) ) ;
    nor_HPC2 SboxInst_U289 ( .a ({new_AGEMA_signal_2593, y0[38]}), .b ({new_AGEMA_signal_2958, SboxInst_n225}), .clk (clk), .r (Fresh[159]), .c ({new_AGEMA_signal_3142, z4[38]}) ) ;
    nor_HPC2 SboxInst_U288 ( .a ({new_AGEMA_signal_2591, y0[39]}), .b ({new_AGEMA_signal_2916, SboxInst_n224}), .clk (clk), .r (Fresh[160]), .c ({new_AGEMA_signal_3143, z4[39]}) ) ;
    nor_HPC2 SboxInst_U287 ( .a ({new_AGEMA_signal_2589, y0[3]}), .b ({new_AGEMA_signal_2904, SboxInst_n223}), .clk (clk), .r (Fresh[161]), .c ({new_AGEMA_signal_3144, z4[3]}) ) ;
    nor_HPC2 SboxInst_U286 ( .a ({new_AGEMA_signal_2587, y0[40]}), .b ({new_AGEMA_signal_2914, SboxInst_n222}), .clk (clk), .r (Fresh[162]), .c ({new_AGEMA_signal_3145, z4[40]}) ) ;
    nor_HPC2 SboxInst_U285 ( .a ({new_AGEMA_signal_2585, y0[41]}), .b ({new_AGEMA_signal_2913, SboxInst_n221}), .clk (clk), .r (Fresh[163]), .c ({new_AGEMA_signal_3146, z4[41]}) ) ;
    nor_HPC2 SboxInst_U284 ( .a ({new_AGEMA_signal_2583, y0[42]}), .b ({new_AGEMA_signal_2910, SboxInst_n220}), .clk (clk), .r (Fresh[164]), .c ({new_AGEMA_signal_3147, z4[42]}) ) ;
    nor_HPC2 SboxInst_U283 ( .a ({new_AGEMA_signal_2581, y0[43]}), .b ({new_AGEMA_signal_2908, SboxInst_n219}), .clk (clk), .r (Fresh[165]), .c ({new_AGEMA_signal_3148, z4[43]}) ) ;
    nor_HPC2 SboxInst_U282 ( .a ({new_AGEMA_signal_2579, y0[44]}), .b ({new_AGEMA_signal_2905, SboxInst_n218}), .clk (clk), .r (Fresh[166]), .c ({new_AGEMA_signal_3149, z4[44]}) ) ;
    nor_HPC2 SboxInst_U281 ( .a ({new_AGEMA_signal_2577, y0[45]}), .b ({new_AGEMA_signal_2902, SboxInst_n217}), .clk (clk), .r (Fresh[167]), .c ({new_AGEMA_signal_3150, z4[45]}) ) ;
    nor_HPC2 SboxInst_U280 ( .a ({new_AGEMA_signal_2575, y0[46]}), .b ({new_AGEMA_signal_2897, SboxInst_n216}), .clk (clk), .r (Fresh[168]), .c ({new_AGEMA_signal_3151, z4[46]}) ) ;
    nor_HPC2 SboxInst_U279 ( .a ({new_AGEMA_signal_2573, y0[47]}), .b ({new_AGEMA_signal_2933, SboxInst_n215}), .clk (clk), .r (Fresh[169]), .c ({new_AGEMA_signal_3152, z4[47]}) ) ;
    nor_HPC2 SboxInst_U278 ( .a ({new_AGEMA_signal_2571, y0[48]}), .b ({new_AGEMA_signal_2932, SboxInst_n214}), .clk (clk), .r (Fresh[170]), .c ({new_AGEMA_signal_3153, z4[48]}) ) ;
    nor_HPC2 SboxInst_U277 ( .a ({new_AGEMA_signal_2569, y0[49]}), .b ({new_AGEMA_signal_2931, SboxInst_n213}), .clk (clk), .r (Fresh[171]), .c ({new_AGEMA_signal_3154, z4[49]}) ) ;
    nor_HPC2 SboxInst_U276 ( .a ({new_AGEMA_signal_2567, y0[4]}), .b ({new_AGEMA_signal_2900, SboxInst_n212}), .clk (clk), .r (Fresh[172]), .c ({new_AGEMA_signal_3155, z4[4]}) ) ;
    nor_HPC2 SboxInst_U275 ( .a ({new_AGEMA_signal_2565, y0[50]}), .b ({new_AGEMA_signal_2930, SboxInst_n211}), .clk (clk), .r (Fresh[173]), .c ({new_AGEMA_signal_3156, z4[50]}) ) ;
    nor_HPC2 SboxInst_U274 ( .a ({new_AGEMA_signal_2563, y0[51]}), .b ({new_AGEMA_signal_2928, SboxInst_n210}), .clk (clk), .r (Fresh[174]), .c ({new_AGEMA_signal_3157, z4[51]}) ) ;
    nor_HPC2 SboxInst_U273 ( .a ({new_AGEMA_signal_2561, y0[52]}), .b ({new_AGEMA_signal_2926, SboxInst_n209}), .clk (clk), .r (Fresh[175]), .c ({new_AGEMA_signal_3158, z4[52]}) ) ;
    nor_HPC2 SboxInst_U272 ( .a ({new_AGEMA_signal_2559, y0[53]}), .b ({new_AGEMA_signal_2923, SboxInst_n208}), .clk (clk), .r (Fresh[176]), .c ({new_AGEMA_signal_3159, z4[53]}) ) ;
    nor_HPC2 SboxInst_U271 ( .a ({new_AGEMA_signal_2557, y0[54]}), .b ({new_AGEMA_signal_2920, SboxInst_n207}), .clk (clk), .r (Fresh[177]), .c ({new_AGEMA_signal_3160, z4[54]}) ) ;
    nor_HPC2 SboxInst_U270 ( .a ({new_AGEMA_signal_2555, y0[55]}), .b ({new_AGEMA_signal_2947, SboxInst_n206}), .clk (clk), .r (Fresh[178]), .c ({new_AGEMA_signal_3161, z4[55]}) ) ;
    nor_HPC2 SboxInst_U269 ( .a ({new_AGEMA_signal_2553, y0[56]}), .b ({new_AGEMA_signal_2946, SboxInst_n205}), .clk (clk), .r (Fresh[179]), .c ({new_AGEMA_signal_3162, z4[56]}) ) ;
    nor_HPC2 SboxInst_U268 ( .a ({new_AGEMA_signal_2551, y0[57]}), .b ({new_AGEMA_signal_2945, SboxInst_n204}), .clk (clk), .r (Fresh[180]), .c ({new_AGEMA_signal_3163, z4[57]}) ) ;
    nor_HPC2 SboxInst_U267 ( .a ({new_AGEMA_signal_2549, y0[58]}), .b ({new_AGEMA_signal_2943, SboxInst_n203}), .clk (clk), .r (Fresh[181]), .c ({new_AGEMA_signal_3164, z4[58]}) ) ;
    nor_HPC2 SboxInst_U266 ( .a ({new_AGEMA_signal_2547, y0[59]}), .b ({new_AGEMA_signal_2941, SboxInst_n202}), .clk (clk), .r (Fresh[182]), .c ({new_AGEMA_signal_3165, z4[59]}) ) ;
    nor_HPC2 SboxInst_U265 ( .a ({new_AGEMA_signal_2545, y0[5]}), .b ({new_AGEMA_signal_2907, SboxInst_n201}), .clk (clk), .r (Fresh[183]), .c ({new_AGEMA_signal_3166, z4[5]}) ) ;
    nor_HPC2 SboxInst_U264 ( .a ({new_AGEMA_signal_2543, y0[60]}), .b ({new_AGEMA_signal_2938, SboxInst_n200}), .clk (clk), .r (Fresh[184]), .c ({new_AGEMA_signal_3167, z4[60]}) ) ;
    nor_HPC2 SboxInst_U263 ( .a ({new_AGEMA_signal_2541, y0[61]}), .b ({new_AGEMA_signal_2917, SboxInst_n199}), .clk (clk), .r (Fresh[185]), .c ({new_AGEMA_signal_3168, z4[61]}) ) ;
    nor_HPC2 SboxInst_U262 ( .a ({new_AGEMA_signal_2539, y0[62]}), .b ({new_AGEMA_signal_2915, SboxInst_n198}), .clk (clk), .r (Fresh[186]), .c ({new_AGEMA_signal_3169, z4[62]}) ) ;
    nor_HPC2 SboxInst_U261 ( .a ({new_AGEMA_signal_2537, y0[63]}), .b ({new_AGEMA_signal_2912, SboxInst_n197}), .clk (clk), .r (Fresh[187]), .c ({new_AGEMA_signal_3170, z4[63]}) ) ;
    nor_HPC2 SboxInst_U260 ( .a ({new_AGEMA_signal_2535, y0[6]}), .b ({new_AGEMA_signal_2901, SboxInst_n196}), .clk (clk), .r (Fresh[188]), .c ({new_AGEMA_signal_3171, z4[6]}) ) ;
    nor_HPC2 SboxInst_U259 ( .a ({new_AGEMA_signal_2533, y0[7]}), .b ({new_AGEMA_signal_2899, SboxInst_n195}), .clk (clk), .r (Fresh[189]), .c ({new_AGEMA_signal_3172, z4[7]}) ) ;
    nor_HPC2 SboxInst_U258 ( .a ({new_AGEMA_signal_2531, y0[8]}), .b ({new_AGEMA_signal_2929, SboxInst_n194}), .clk (clk), .r (Fresh[190]), .c ({new_AGEMA_signal_3173, z4[8]}) ) ;
    nor_HPC2 SboxInst_U257 ( .a ({new_AGEMA_signal_2529, y0[9]}), .b ({new_AGEMA_signal_2927, SboxInst_n193}), .clk (clk), .r (Fresh[191]), .c ({new_AGEMA_signal_3174, z4[9]}) ) ;
    and_HPC2 SboxInst_U256 ( .a ({new_AGEMA_signal_2859, SboxInst_n345}), .b ({new_AGEMA_signal_2410, y4[45]}), .clk (clk), .r (Fresh[192]), .c ({new_AGEMA_signal_3175, z2[45]}) ) ;
    and_HPC2 SboxInst_U254 ( .a ({new_AGEMA_signal_2860, SboxInst_n352}), .b ({new_AGEMA_signal_2431, y4[39]}), .clk (clk), .r (Fresh[193]), .c ({new_AGEMA_signal_3176, z2[39]}) ) ;
    and_HPC2 SboxInst_U252 ( .a ({new_AGEMA_signal_2861, SboxInst_n350}), .b ({new_AGEMA_signal_2425, y4[40]}), .clk (clk), .r (Fresh[194]), .c ({new_AGEMA_signal_3177, z2[40]}) ) ;
    and_HPC2 SboxInst_U250 ( .a ({new_AGEMA_signal_2862, SboxInst_n346}), .b ({new_AGEMA_signal_2413, y4[44]}), .clk (clk), .r (Fresh[195]), .c ({new_AGEMA_signal_3178, z2[44]}) ) ;
    and_HPC2 SboxInst_U248 ( .a ({new_AGEMA_signal_2863, SboxInst_n353}), .b ({new_AGEMA_signal_2434, y4[38]}), .clk (clk), .r (Fresh[196]), .c ({new_AGEMA_signal_3179, z2[38]}) ) ;
    and_HPC2 SboxInst_U246 ( .a ({new_AGEMA_signal_2864, SboxInst_n347}), .b ({new_AGEMA_signal_2416, y4[43]}), .clk (clk), .r (Fresh[197]), .c ({new_AGEMA_signal_3180, z2[43]}) ) ;
    and_HPC2 SboxInst_U244 ( .a ({new_AGEMA_signal_2865, SboxInst_n354}), .b ({new_AGEMA_signal_2437, y4[37]}), .clk (clk), .r (Fresh[198]), .c ({new_AGEMA_signal_3181, z2[37]}) ) ;
    and_HPC2 SboxInst_U242 ( .a ({new_AGEMA_signal_2866, SboxInst_n348}), .b ({new_AGEMA_signal_2419, y4[42]}), .clk (clk), .r (Fresh[199]), .c ({new_AGEMA_signal_3182, z2[42]}) ) ;
    and_HPC2 SboxInst_U240 ( .a ({new_AGEMA_signal_2867, SboxInst_n355}), .b ({new_AGEMA_signal_2440, y4[36]}), .clk (clk), .r (Fresh[200]), .c ({new_AGEMA_signal_3183, z2[36]}) ) ;
    and_HPC2 SboxInst_U238 ( .a ({new_AGEMA_signal_2868, SboxInst_n349}), .b ({new_AGEMA_signal_2422, y4[41]}), .clk (clk), .r (Fresh[201]), .c ({new_AGEMA_signal_3184, z2[41]}) ) ;
    and_HPC2 SboxInst_U236 ( .a ({new_AGEMA_signal_2869, SboxInst_n356}), .b ({new_AGEMA_signal_2443, y4[35]}), .clk (clk), .r (Fresh[202]), .c ({new_AGEMA_signal_3185, z2[35]}) ) ;
    and_HPC2 SboxInst_U234 ( .a ({new_AGEMA_signal_2870, SboxInst_n357}), .b ({new_AGEMA_signal_2446, y4[34]}), .clk (clk), .r (Fresh[203]), .c ({new_AGEMA_signal_3186, z2[34]}) ) ;
    and_HPC2 SboxInst_U232 ( .a ({new_AGEMA_signal_2871, SboxInst_n358}), .b ({new_AGEMA_signal_2449, y4[33]}), .clk (clk), .r (Fresh[204]), .c ({new_AGEMA_signal_3187, z2[33]}) ) ;
    and_HPC2 SboxInst_U230 ( .a ({new_AGEMA_signal_2872, SboxInst_n359}), .b ({new_AGEMA_signal_2452, y4[32]}), .clk (clk), .r (Fresh[205]), .c ({new_AGEMA_signal_3188, z2[32]}) ) ;
    and_HPC2 SboxInst_U228 ( .a ({new_AGEMA_signal_2873, SboxInst_n342}), .b ({new_AGEMA_signal_2401, y4[48]}), .clk (clk), .r (Fresh[206]), .c ({new_AGEMA_signal_3189, z2[48]}) ) ;
    and_HPC2 SboxInst_U226 ( .a ({new_AGEMA_signal_2874, SboxInst_n336}), .b ({new_AGEMA_signal_2383, y4[53]}), .clk (clk), .r (Fresh[207]), .c ({new_AGEMA_signal_3190, z2[53]}) ) ;
    and_HPC2 SboxInst_U224 ( .a ({new_AGEMA_signal_2875, SboxInst_n343}), .b ({new_AGEMA_signal_2404, y4[47]}), .clk (clk), .r (Fresh[208]), .c ({new_AGEMA_signal_3191, z2[47]}) ) ;
    and_HPC2 SboxInst_U222 ( .a ({new_AGEMA_signal_2876, SboxInst_n337}), .b ({new_AGEMA_signal_2386, y4[52]}), .clk (clk), .r (Fresh[209]), .c ({new_AGEMA_signal_3192, z2[52]}) ) ;
    and_HPC2 SboxInst_U220 ( .a ({new_AGEMA_signal_2877, SboxInst_n344}), .b ({new_AGEMA_signal_2407, y4[46]}), .clk (clk), .r (Fresh[210]), .c ({new_AGEMA_signal_3193, z2[46]}) ) ;
    and_HPC2 SboxInst_U218 ( .a ({new_AGEMA_signal_2878, SboxInst_n338}), .b ({new_AGEMA_signal_2389, y4[51]}), .clk (clk), .r (Fresh[211]), .c ({new_AGEMA_signal_3194, z2[51]}) ) ;
    and_HPC2 SboxInst_U216 ( .a ({new_AGEMA_signal_2879, SboxInst_n339}), .b ({new_AGEMA_signal_2392, y4[50]}), .clk (clk), .r (Fresh[212]), .c ({new_AGEMA_signal_3195, z2[50]}) ) ;
    and_HPC2 SboxInst_U214 ( .a ({new_AGEMA_signal_2880, SboxInst_n341}), .b ({new_AGEMA_signal_2398, y4[49]}), .clk (clk), .r (Fresh[213]), .c ({new_AGEMA_signal_3196, z2[49]}) ) ;
    and_HPC2 SboxInst_U212 ( .a ({new_AGEMA_signal_2881, SboxInst_n334}), .b ({new_AGEMA_signal_2377, y4[55]}), .clk (clk), .r (Fresh[214]), .c ({new_AGEMA_signal_3197, z2[55]}) ) ;
    and_HPC2 SboxInst_U210 ( .a ({new_AGEMA_signal_2882, SboxInst_n327}), .b ({new_AGEMA_signal_2356, y4[61]}), .clk (clk), .r (Fresh[215]), .c ({new_AGEMA_signal_3198, z2[61]}) ) ;
    and_HPC2 SboxInst_U208 ( .a ({new_AGEMA_signal_2883, SboxInst_n333}), .b ({new_AGEMA_signal_2374, y4[56]}), .clk (clk), .r (Fresh[216]), .c ({new_AGEMA_signal_3199, z2[56]}) ) ;
    and_HPC2 SboxInst_U206 ( .a ({new_AGEMA_signal_2884, SboxInst_n335}), .b ({new_AGEMA_signal_2380, y4[54]}), .clk (clk), .r (Fresh[217]), .c ({new_AGEMA_signal_3200, z2[54]}) ) ;
    and_HPC2 SboxInst_U204 ( .a ({new_AGEMA_signal_2885, SboxInst_n328}), .b ({new_AGEMA_signal_2359, y4[60]}), .clk (clk), .r (Fresh[218]), .c ({new_AGEMA_signal_3201, z2[60]}) ) ;
    and_HPC2 SboxInst_U202 ( .a ({new_AGEMA_signal_2886, SboxInst_n330}), .b ({new_AGEMA_signal_2365, y4[59]}), .clk (clk), .r (Fresh[219]), .c ({new_AGEMA_signal_3202, z2[59]}) ) ;
    and_HPC2 SboxInst_U200 ( .a ({new_AGEMA_signal_2887, SboxInst_n331}), .b ({new_AGEMA_signal_2368, y4[58]}), .clk (clk), .r (Fresh[220]), .c ({new_AGEMA_signal_3203, z2[58]}) ) ;
    and_HPC2 SboxInst_U198 ( .a ({new_AGEMA_signal_2888, SboxInst_n332}), .b ({new_AGEMA_signal_2371, y4[57]}), .clk (clk), .r (Fresh[221]), .c ({new_AGEMA_signal_3204, z2[57]}) ) ;
    and_HPC2 SboxInst_U196 ( .a ({new_AGEMA_signal_2889, SboxInst_n325}), .b ({new_AGEMA_signal_2350, y4[63]}), .clk (clk), .r (Fresh[222]), .c ({new_AGEMA_signal_3205, z2[63]}) ) ;
    and_HPC2 SboxInst_U194 ( .a ({new_AGEMA_signal_2890, SboxInst_n384}), .b ({new_AGEMA_signal_2527, y4[0]}), .clk (clk), .r (Fresh[223]), .c ({new_AGEMA_signal_3206, z2[0]}) ) ;
    and_HPC2 SboxInst_U192 ( .a ({new_AGEMA_signal_2891, SboxInst_n329}), .b ({new_AGEMA_signal_2362, y4[5]}), .clk (clk), .r (Fresh[224]), .c ({new_AGEMA_signal_3207, z2[5]}) ) ;
    and_HPC2 SboxInst_U190 ( .a ({new_AGEMA_signal_2892, SboxInst_n340}), .b ({new_AGEMA_signal_2395, y4[4]}), .clk (clk), .r (Fresh[225]), .c ({new_AGEMA_signal_3208, z2[4]}) ) ;
    and_HPC2 SboxInst_U188 ( .a ({new_AGEMA_signal_2893, SboxInst_n326}), .b ({new_AGEMA_signal_2353, y4[62]}), .clk (clk), .r (Fresh[226]), .c ({new_AGEMA_signal_3209, z2[62]}) ) ;
    and_HPC2 SboxInst_U186 ( .a ({new_AGEMA_signal_2894, SboxInst_n351}), .b ({new_AGEMA_signal_2428, y4[3]}), .clk (clk), .r (Fresh[227]), .c ({new_AGEMA_signal_3210, z2[3]}) ) ;
    and_HPC2 SboxInst_U184 ( .a ({new_AGEMA_signal_2895, SboxInst_n362}), .b ({new_AGEMA_signal_2461, y4[2]}), .clk (clk), .r (Fresh[228]), .c ({new_AGEMA_signal_3211, z2[2]}) ) ;
    and_HPC2 SboxInst_U182 ( .a ({new_AGEMA_signal_2896, SboxInst_n373}), .b ({new_AGEMA_signal_2494, y4[1]}), .clk (clk), .r (Fresh[229]), .c ({new_AGEMA_signal_3212, z2[1]}) ) ;
    and_HPC2 SboxInst_U180 ( .a ({new_AGEMA_signal_2793, n3253}), .b ({new_AGEMA_signal_2897, SboxInst_n216}), .clk (clk), .r (Fresh[230]), .c ({new_AGEMA_signal_3213, z0[46]}) ) ;
    and_HPC2 SboxInst_U178 ( .a ({new_AGEMA_signal_4433, n3239}), .b ({new_AGEMA_signal_2899, SboxInst_n195}), .clk (clk), .r (Fresh[231]), .c ({new_AGEMA_signal_4579, z0[7]}) ) ;
    and_HPC2 SboxInst_U176 ( .a ({new_AGEMA_signal_2990, n3232}), .b ({new_AGEMA_signal_2900, SboxInst_n212}), .clk (clk), .r (Fresh[232]), .c ({new_AGEMA_signal_3583, z0[4]}) ) ;
    and_HPC2 SboxInst_U174 ( .a ({new_AGEMA_signal_3826, n3230}), .b ({new_AGEMA_signal_2901, SboxInst_n196}), .clk (clk), .r (Fresh[233]), .c ({new_AGEMA_signal_4202, z0[6]}) ) ;
    and_HPC2 SboxInst_U172 ( .a ({new_AGEMA_signal_2790, n3254}), .b ({new_AGEMA_signal_2902, SboxInst_n217}), .clk (clk), .r (Fresh[234]), .c ({new_AGEMA_signal_3214, z0[45]}) ) ;
    and_HPC2 SboxInst_U170 ( .a ({new_AGEMA_signal_4432, n3233}), .b ({new_AGEMA_signal_2904, SboxInst_n223}), .clk (clk), .r (Fresh[235]), .c ({new_AGEMA_signal_4580, z0[3]}) ) ;
    and_HPC2 SboxInst_U168 ( .a ({new_AGEMA_signal_2788, n3255}), .b ({new_AGEMA_signal_2905, SboxInst_n218}), .clk (clk), .r (Fresh[236]), .c ({new_AGEMA_signal_3215, z0[44]}) ) ;
    and_HPC2 SboxInst_U166 ( .a ({new_AGEMA_signal_3824, n3287}), .b ({new_AGEMA_signal_2906, SboxInst_n234}), .clk (clk), .r (Fresh[237]), .c ({new_AGEMA_signal_4203, z0[2]}) ) ;
    and_HPC2 SboxInst_U164 ( .a ({new_AGEMA_signal_3515, n3231}), .b ({new_AGEMA_signal_2907, SboxInst_n201}), .clk (clk), .r (Fresh[238]), .c ({new_AGEMA_signal_3889, z0[5]}) ) ;
    and_HPC2 SboxInst_U162 ( .a ({new_AGEMA_signal_2786, n3256}), .b ({new_AGEMA_signal_2908, SboxInst_n219}), .clk (clk), .r (Fresh[239]), .c ({new_AGEMA_signal_3216, z0[43]}) ) ;
    and_HPC2 SboxInst_U160 ( .a ({new_AGEMA_signal_3513, y2[1]}), .b ({new_AGEMA_signal_2909, SboxInst_n245}), .clk (clk), .r (Fresh[240]), .c ({new_AGEMA_signal_3890, z0[1]}) ) ;
    and_HPC2 SboxInst_U158 ( .a ({new_AGEMA_signal_2783, n3257}), .b ({new_AGEMA_signal_2910, SboxInst_n220}), .clk (clk), .r (Fresh[241]), .c ({new_AGEMA_signal_3217, z0[42]}) ) ;
    and_HPC2 SboxInst_U156 ( .a ({new_AGEMA_signal_2989, y2[0]}), .b ({new_AGEMA_signal_2911, SboxInst_n256}), .clk (clk), .r (Fresh[242]), .c ({new_AGEMA_signal_3584, z0[0]}) ) ;
    and_HPC2 SboxInst_U154 ( .a ({new_AGEMA_signal_2846, n3234}), .b ({new_AGEMA_signal_2912, SboxInst_n197}), .clk (clk), .r (Fresh[243]), .c ({new_AGEMA_signal_3218, z0[63]}) ) ;
    and_HPC2 SboxInst_U152 ( .a ({new_AGEMA_signal_2780, n3258}), .b ({new_AGEMA_signal_2913, SboxInst_n221}), .clk (clk), .r (Fresh[244]), .c ({new_AGEMA_signal_3219, z0[41]}) ) ;
    and_HPC2 SboxInst_U150 ( .a ({new_AGEMA_signal_2778, n3259}), .b ({new_AGEMA_signal_2914, SboxInst_n222}), .clk (clk), .r (Fresh[245]), .c ({new_AGEMA_signal_3220, z0[40]}) ) ;
    and_HPC2 SboxInst_U148 ( .a ({new_AGEMA_signal_2840, n3235}), .b ({new_AGEMA_signal_2915, SboxInst_n198}), .clk (clk), .r (Fresh[246]), .c ({new_AGEMA_signal_3221, z0[62]}) ) ;
    and_HPC2 SboxInst_U146 ( .a ({new_AGEMA_signal_2775, n3260}), .b ({new_AGEMA_signal_2916, SboxInst_n224}), .clk (clk), .r (Fresh[247]), .c ({new_AGEMA_signal_3222, z0[39]}) ) ;
    and_HPC2 SboxInst_U144 ( .a ({new_AGEMA_signal_2837, n3236}), .b ({new_AGEMA_signal_2917, SboxInst_n199}), .clk (clk), .r (Fresh[248]), .c ({new_AGEMA_signal_3223, z0[61]}) ) ;
    and_HPC2 SboxInst_U142 ( .a ({new_AGEMA_signal_2742, n3284}), .b ({new_AGEMA_signal_2918, SboxInst_n250}), .clk (clk), .r (Fresh[249]), .c ({new_AGEMA_signal_3224, z0[15]}) ) ;
    and_HPC2 SboxInst_U140 ( .a ({new_AGEMA_signal_2717, n3288}), .b ({new_AGEMA_signal_2919, SboxInst_n253}), .clk (clk), .r (Fresh[250]), .c ({new_AGEMA_signal_3225, z0[12]}) ) ;
    and_HPC2 SboxInst_U138 ( .a ({new_AGEMA_signal_2813, n3245}), .b ({new_AGEMA_signal_2920, SboxInst_n207}), .clk (clk), .r (Fresh[251]), .c ({new_AGEMA_signal_3226, z0[54]}) ) ;
    and_HPC2 SboxInst_U136 ( .a ({new_AGEMA_signal_2709, n3289}), .b ({new_AGEMA_signal_2921, SboxInst_n254}), .clk (clk), .r (Fresh[252]), .c ({new_AGEMA_signal_3227, z0[11]}) ) ;
    and_HPC2 SboxInst_U134 ( .a ({new_AGEMA_signal_2733, n3285}), .b ({new_AGEMA_signal_2922, SboxInst_n251}), .clk (clk), .r (Fresh[253]), .c ({new_AGEMA_signal_3228, z0[14]}) ) ;
    and_HPC2 SboxInst_U132 ( .a ({new_AGEMA_signal_2810, n3246}), .b ({new_AGEMA_signal_2923, SboxInst_n208}), .clk (clk), .r (Fresh[254]), .c ({new_AGEMA_signal_3229, z0[53]}) ) ;
    and_HPC2 SboxInst_U130 ( .a ({new_AGEMA_signal_2704, n3290}), .b ({new_AGEMA_signal_2924, SboxInst_n255}), .clk (clk), .r (Fresh[255]), .c ({new_AGEMA_signal_3230, z0[10]}) ) ;
    and_HPC2 SboxInst_U128 ( .a ({new_AGEMA_signal_2727, n3286}), .b ({new_AGEMA_signal_2925, SboxInst_n252}), .clk (clk), .r (Fresh[256]), .c ({new_AGEMA_signal_3231, z0[13]}) ) ;
    and_HPC2 SboxInst_U126 ( .a ({new_AGEMA_signal_2807, n3247}), .b ({new_AGEMA_signal_2926, SboxInst_n209}), .clk (clk), .r (Fresh[257]), .c ({new_AGEMA_signal_3232, z0[52]}) ) ;
    and_HPC2 SboxInst_U124 ( .a ({new_AGEMA_signal_2692, n3291}), .b ({new_AGEMA_signal_2927, SboxInst_n193}), .clk (clk), .r (Fresh[258]), .c ({new_AGEMA_signal_3233, z0[9]}) ) ;
    and_HPC2 SboxInst_U122 ( .a ({new_AGEMA_signal_2805, n3248}), .b ({new_AGEMA_signal_2928, SboxInst_n210}), .clk (clk), .r (Fresh[259]), .c ({new_AGEMA_signal_3234, z0[51]}) ) ;
    and_HPC2 SboxInst_U120 ( .a ({new_AGEMA_signal_2834, n3237}), .b ({new_AGEMA_signal_2929, SboxInst_n194}), .clk (clk), .r (Fresh[260]), .c ({new_AGEMA_signal_3235, z0[8]}) ) ;
    and_HPC2 SboxInst_U118 ( .a ({new_AGEMA_signal_2803, n3249}), .b ({new_AGEMA_signal_2930, SboxInst_n211}), .clk (clk), .r (Fresh[261]), .c ({new_AGEMA_signal_3236, z0[50]}) ) ;
    and_HPC2 SboxInst_U116 ( .a ({new_AGEMA_signal_2800, n3250}), .b ({new_AGEMA_signal_2931, SboxInst_n213}), .clk (clk), .r (Fresh[262]), .c ({new_AGEMA_signal_3237, z0[49]}) ) ;
    and_HPC2 SboxInst_U114 ( .a ({new_AGEMA_signal_2797, n3251}), .b ({new_AGEMA_signal_2932, SboxInst_n214}), .clk (clk), .r (Fresh[263]), .c ({new_AGEMA_signal_3238, z0[48]}) ) ;
    and_HPC2 SboxInst_U112 ( .a ({new_AGEMA_signal_2795, n3252}), .b ({new_AGEMA_signal_2933, SboxInst_n215}), .clk (clk), .r (Fresh[264]), .c ({new_AGEMA_signal_3239, z0[47]}) ) ;
    and_HPC2 SboxInst_U110 ( .a ({new_AGEMA_signal_2701, n3279}), .b ({new_AGEMA_signal_2934, SboxInst_n244}), .clk (clk), .r (Fresh[265]), .c ({new_AGEMA_signal_3240, z0[20]}) ) ;
    and_HPC2 SboxInst_U108 ( .a ({new_AGEMA_signal_2724, n3276}), .b ({new_AGEMA_signal_2935, SboxInst_n241}), .clk (clk), .r (Fresh[266]), .c ({new_AGEMA_signal_3241, z0[23]}) ) ;
    and_HPC2 SboxInst_U106 ( .a ({new_AGEMA_signal_2695, n3280}), .b ({new_AGEMA_signal_2936, SboxInst_n246}), .clk (clk), .r (Fresh[267]), .c ({new_AGEMA_signal_3242, z0[19]}) ) ;
    and_HPC2 SboxInst_U104 ( .a ({new_AGEMA_signal_2719, n3277}), .b ({new_AGEMA_signal_2937, SboxInst_n242}), .clk (clk), .r (Fresh[268]), .c ({new_AGEMA_signal_3243, z0[22]}) ) ;
    and_HPC2 SboxInst_U102 ( .a ({new_AGEMA_signal_2828, n3238}), .b ({new_AGEMA_signal_2938, SboxInst_n200}), .clk (clk), .r (Fresh[269]), .c ({new_AGEMA_signal_3244, z0[60]}) ) ;
    and_HPC2 SboxInst_U100 ( .a ({new_AGEMA_signal_2712, n3278}), .b ({new_AGEMA_signal_2939, SboxInst_n243}), .clk (clk), .r (Fresh[270]), .c ({new_AGEMA_signal_3245, z0[21]}) ) ;
    and_HPC2 SboxInst_U98 ( .a ({new_AGEMA_signal_2760, n3281}), .b ({new_AGEMA_signal_2940, SboxInst_n247}), .clk (clk), .r (Fresh[271]), .c ({new_AGEMA_signal_3246, z0[18]}) ) ;
    and_HPC2 SboxInst_U96 ( .a ({new_AGEMA_signal_2825, n3240}), .b ({new_AGEMA_signal_2941, SboxInst_n202}), .clk (clk), .r (Fresh[272]), .c ({new_AGEMA_signal_3247, z0[59]}) ) ;
    and_HPC2 SboxInst_U94 ( .a ({new_AGEMA_signal_2755, n3282}), .b ({new_AGEMA_signal_2942, SboxInst_n248}), .clk (clk), .r (Fresh[273]), .c ({new_AGEMA_signal_3248, z0[17]}) ) ;
    and_HPC2 SboxInst_U92 ( .a ({new_AGEMA_signal_2823, n3241}), .b ({new_AGEMA_signal_2943, SboxInst_n203}), .clk (clk), .r (Fresh[274]), .c ({new_AGEMA_signal_3249, z0[58]}) ) ;
    and_HPC2 SboxInst_U90 ( .a ({new_AGEMA_signal_2750, n3283}), .b ({new_AGEMA_signal_2944, SboxInst_n249}), .clk (clk), .r (Fresh[275]), .c ({new_AGEMA_signal_3250, z0[16]}) ) ;
    and_HPC2 SboxInst_U88 ( .a ({new_AGEMA_signal_2821, n3242}), .b ({new_AGEMA_signal_2945, SboxInst_n204}), .clk (clk), .r (Fresh[276]), .c ({new_AGEMA_signal_3251, z0[57]}) ) ;
    and_HPC2 SboxInst_U86 ( .a ({new_AGEMA_signal_2819, n3243}), .b ({new_AGEMA_signal_2946, SboxInst_n205}), .clk (clk), .r (Fresh[277]), .c ({new_AGEMA_signal_3252, z0[56]}) ) ;
    and_HPC2 SboxInst_U84 ( .a ({new_AGEMA_signal_2816, n3244}), .b ({new_AGEMA_signal_2947, SboxInst_n206}), .clk (clk), .r (Fresh[278]), .c ({new_AGEMA_signal_3253, z0[55]}) ) ;
    and_HPC2 SboxInst_U82 ( .a ({new_AGEMA_signal_2739, n3268}), .b ({new_AGEMA_signal_2948, SboxInst_n232}), .clk (clk), .r (Fresh[279]), .c ({new_AGEMA_signal_3254, z0[31]}) ) ;
    and_HPC2 SboxInst_U80 ( .a ({new_AGEMA_signal_2714, n3271}), .b ({new_AGEMA_signal_2949, SboxInst_n236}), .clk (clk), .r (Fresh[280]), .c ({new_AGEMA_signal_3255, z0[28]}) ) ;
    and_HPC2 SboxInst_U78 ( .a ({new_AGEMA_signal_2730, n3269}), .b ({new_AGEMA_signal_2950, SboxInst_n233}), .clk (clk), .r (Fresh[281]), .c ({new_AGEMA_signal_3256, z0[30]}) ) ;
    and_HPC2 SboxInst_U76 ( .a ({new_AGEMA_signal_2707, n3272}), .b ({new_AGEMA_signal_2951, SboxInst_n237}), .clk (clk), .r (Fresh[282]), .c ({new_AGEMA_signal_3257, z0[27]}) ) ;
    and_HPC2 SboxInst_U74 ( .a ({new_AGEMA_signal_2698, n3273}), .b ({new_AGEMA_signal_2952, SboxInst_n238}), .clk (clk), .r (Fresh[283]), .c ({new_AGEMA_signal_3258, z0[26]}) ) ;
    and_HPC2 SboxInst_U72 ( .a ({new_AGEMA_signal_2721, n3270}), .b ({new_AGEMA_signal_2953, SboxInst_n235}), .clk (clk), .r (Fresh[284]), .c ({new_AGEMA_signal_3259, z0[29]}) ) ;
    and_HPC2 SboxInst_U70 ( .a ({new_AGEMA_signal_2744, n3274}), .b ({new_AGEMA_signal_2954, SboxInst_n239}), .clk (clk), .r (Fresh[285]), .c ({new_AGEMA_signal_3260, z0[25]}) ) ;
    and_HPC2 SboxInst_U68 ( .a ({new_AGEMA_signal_2736, n3275}), .b ({new_AGEMA_signal_2955, SboxInst_n240}), .clk (clk), .r (Fresh[286]), .c ({new_AGEMA_signal_3261, z0[24]}) ) ;
    and_HPC2 SboxInst_U66 ( .a ({new_AGEMA_signal_2766, n3263}), .b ({new_AGEMA_signal_2956, SboxInst_n227}), .clk (clk), .r (Fresh[287]), .c ({new_AGEMA_signal_3262, z0[36]}) ) ;
    and_HPC2 SboxInst_U64 ( .a ({new_AGEMA_signal_2763, n3264}), .b ({new_AGEMA_signal_2957, SboxInst_n228}), .clk (clk), .r (Fresh[288]), .c ({new_AGEMA_signal_3263, z0[35]}) ) ;
    and_HPC2 SboxInst_U62 ( .a ({new_AGEMA_signal_2772, n3261}), .b ({new_AGEMA_signal_2958, SboxInst_n225}), .clk (clk), .r (Fresh[289]), .c ({new_AGEMA_signal_3264, z0[38]}) ) ;
    and_HPC2 SboxInst_U60 ( .a ({new_AGEMA_signal_2758, n3265}), .b ({new_AGEMA_signal_2959, SboxInst_n229}), .clk (clk), .r (Fresh[290]), .c ({new_AGEMA_signal_3265, z0[34]}) ) ;
    and_HPC2 SboxInst_U58 ( .a ({new_AGEMA_signal_2769, n3262}), .b ({new_AGEMA_signal_2960, SboxInst_n226}), .clk (clk), .r (Fresh[291]), .c ({new_AGEMA_signal_3266, z0[37]}) ) ;
    and_HPC2 SboxInst_U56 ( .a ({new_AGEMA_signal_2753, n3266}), .b ({new_AGEMA_signal_2961, SboxInst_n230}), .clk (clk), .r (Fresh[292]), .c ({new_AGEMA_signal_3267, z0[33]}) ) ;
    and_HPC2 SboxInst_U54 ( .a ({new_AGEMA_signal_2747, n3267}), .b ({new_AGEMA_signal_2962, SboxInst_n231}), .clk (clk), .r (Fresh[293]), .c ({new_AGEMA_signal_3268, z0[32]}) ) ;
    and_HPC2 SboxInst_U52 ( .a ({new_AGEMA_signal_2963, SboxInst_n323}), .b ({new_AGEMA_signal_2344, y4[7]}), .clk (clk), .r (Fresh[294]), .c ({new_AGEMA_signal_3269, z2[7]}) ) ;
    and_HPC2 SboxInst_U50 ( .a ({new_AGEMA_signal_2964, SboxInst_n376}), .b ({new_AGEMA_signal_2503, y4[17]}), .clk (clk), .r (Fresh[295]), .c ({new_AGEMA_signal_3270, z2[17]}) ) ;
    and_HPC2 SboxInst_U48 ( .a ({new_AGEMA_signal_2965, SboxInst_n368}), .b ({new_AGEMA_signal_2479, y4[24]}), .clk (clk), .r (Fresh[296]), .c ({new_AGEMA_signal_3271, z2[24]}) ) ;
    and_HPC2 SboxInst_U46 ( .a ({new_AGEMA_signal_2966, SboxInst_n324}), .b ({new_AGEMA_signal_2347, y4[6]}), .clk (clk), .r (Fresh[297]), .c ({new_AGEMA_signal_3272, z2[6]}) ) ;
    and_HPC2 SboxInst_U44 ( .a ({new_AGEMA_signal_2967, SboxInst_n369}), .b ({new_AGEMA_signal_2482, y4[23]}), .clk (clk), .r (Fresh[298]), .c ({new_AGEMA_signal_3273, z2[23]}) ) ;
    and_HPC2 SboxInst_U42 ( .a ({new_AGEMA_signal_2968, SboxInst_n377}), .b ({new_AGEMA_signal_2506, y4[16]}), .clk (clk), .r (Fresh[299]), .c ({new_AGEMA_signal_3274, z2[16]}) ) ;
    and_HPC2 SboxInst_U40 ( .a ({new_AGEMA_signal_2969, SboxInst_n370}), .b ({new_AGEMA_signal_2485, y4[22]}), .clk (clk), .r (Fresh[300]), .c ({new_AGEMA_signal_3275, z2[22]}) ) ;
    and_HPC2 SboxInst_U38 ( .a ({new_AGEMA_signal_2970, SboxInst_n378}), .b ({new_AGEMA_signal_2509, y4[15]}), .clk (clk), .r (Fresh[301]), .c ({new_AGEMA_signal_3276, z2[15]}) ) ;
    and_HPC2 SboxInst_U36 ( .a ({new_AGEMA_signal_2971, SboxInst_n379}), .b ({new_AGEMA_signal_2512, y4[14]}), .clk (clk), .r (Fresh[302]), .c ({new_AGEMA_signal_3277, z2[14]}) ) ;
    and_HPC2 SboxInst_U34 ( .a ({new_AGEMA_signal_2972, SboxInst_n371}), .b ({new_AGEMA_signal_2488, y4[21]}), .clk (clk), .r (Fresh[303]), .c ({new_AGEMA_signal_3278, z2[21]}) ) ;
    and_HPC2 SboxInst_U32 ( .a ({new_AGEMA_signal_2973, SboxInst_n372}), .b ({new_AGEMA_signal_2491, y4[20]}), .clk (clk), .r (Fresh[304]), .c ({new_AGEMA_signal_3279, z2[20]}) ) ;
    and_HPC2 SboxInst_U30 ( .a ({new_AGEMA_signal_2974, SboxInst_n380}), .b ({new_AGEMA_signal_2515, y4[13]}), .clk (clk), .r (Fresh[305]), .c ({new_AGEMA_signal_3280, z2[13]}) ) ;
    and_HPC2 SboxInst_U28 ( .a ({new_AGEMA_signal_2975, SboxInst_n381}), .b ({new_AGEMA_signal_2518, y4[12]}), .clk (clk), .r (Fresh[306]), .c ({new_AGEMA_signal_3281, z2[12]}) ) ;
    and_HPC2 SboxInst_U26 ( .a ({new_AGEMA_signal_2976, SboxInst_n374}), .b ({new_AGEMA_signal_2497, y4[19]}), .clk (clk), .r (Fresh[307]), .c ({new_AGEMA_signal_3282, z2[19]}) ) ;
    and_HPC2 SboxInst_U24 ( .a ({new_AGEMA_signal_2977, SboxInst_n382}), .b ({new_AGEMA_signal_2521, y4[11]}), .clk (clk), .r (Fresh[308]), .c ({new_AGEMA_signal_3283, z2[11]}) ) ;
    and_HPC2 SboxInst_U22 ( .a ({new_AGEMA_signal_2978, SboxInst_n375}), .b ({new_AGEMA_signal_2500, y4[18]}), .clk (clk), .r (Fresh[309]), .c ({new_AGEMA_signal_3284, z2[18]}) ) ;
    and_HPC2 SboxInst_U20 ( .a ({new_AGEMA_signal_2979, SboxInst_n383}), .b ({new_AGEMA_signal_2524, y4[10]}), .clk (clk), .r (Fresh[310]), .c ({new_AGEMA_signal_3285, z2[10]}) ) ;
    and_HPC2 SboxInst_U18 ( .a ({new_AGEMA_signal_2980, SboxInst_n367}), .b ({new_AGEMA_signal_2476, y4[25]}), .clk (clk), .r (Fresh[311]), .c ({new_AGEMA_signal_3286, z2[25]}) ) ;
    and_HPC2 SboxInst_U16 ( .a ({new_AGEMA_signal_2981, SboxInst_n360}), .b ({new_AGEMA_signal_2455, y4[31]}), .clk (clk), .r (Fresh[312]), .c ({new_AGEMA_signal_3287, z2[31]}) ) ;
    and_HPC2 SboxInst_U14 ( .a ({new_AGEMA_signal_2982, SboxInst_n361}), .b ({new_AGEMA_signal_2458, y4[30]}), .clk (clk), .r (Fresh[313]), .c ({new_AGEMA_signal_3288, z2[30]}) ) ;
    and_HPC2 SboxInst_U12 ( .a ({new_AGEMA_signal_2983, SboxInst_n363}), .b ({new_AGEMA_signal_2464, y4[29]}), .clk (clk), .r (Fresh[314]), .c ({new_AGEMA_signal_3289, z2[29]}) ) ;
    and_HPC2 SboxInst_U10 ( .a ({new_AGEMA_signal_2984, SboxInst_n364}), .b ({new_AGEMA_signal_2467, y4[28]}), .clk (clk), .r (Fresh[315]), .c ({new_AGEMA_signal_3290, z2[28]}) ) ;
    and_HPC2 SboxInst_U8 ( .a ({new_AGEMA_signal_2985, SboxInst_n365}), .b ({new_AGEMA_signal_2470, y4[27]}), .clk (clk), .r (Fresh[316]), .c ({new_AGEMA_signal_3291, z2[27]}) ) ;
    and_HPC2 SboxInst_U6 ( .a ({new_AGEMA_signal_2986, SboxInst_n321}), .b ({new_AGEMA_signal_2338, y4[9]}), .clk (clk), .r (Fresh[317]), .c ({new_AGEMA_signal_3292, z2[9]}) ) ;
    and_HPC2 SboxInst_U4 ( .a ({new_AGEMA_signal_2987, SboxInst_n366}), .b ({new_AGEMA_signal_2473, y4[26]}), .clk (clk), .r (Fresh[318]), .c ({new_AGEMA_signal_3293, z2[26]}) ) ;
    and_HPC2 SboxInst_U2 ( .a ({new_AGEMA_signal_2988, SboxInst_n322}), .b ({new_AGEMA_signal_2341, y4[8]}), .clk (clk), .r (Fresh[319]), .c ({new_AGEMA_signal_3294, z2[8]}) ) ;

endmodule
