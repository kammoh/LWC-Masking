-- This VHDL was converted from Verilog using the
-- Icarus Verilog VHDL Code Generator 12.0

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Generated from Verilog module Asconp_HPC2_ClockGating_d1 (Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:6)
entity Asconp_HPC2_ClockGating_d1 is
  port (
    clk          : in  std_logic;
    fresh        : in  std_logic_vector(319 downto 0);
    rcon         : in  std_logic_vector(3 downto 0);
    state_in_s0  : in  std_logic_vector(319 downto 0);
    state_in_s1  : in  std_logic_vector(319 downto 0);
    state_out_s0 : out std_logic_vector(319 downto 0);
    state_out_s1 : out std_logic_vector(319 downto 0)
  );
end entity; 

-- Generated from Verilog module Asconp_HPC2_ClockGating_d1 (Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:6)
architecture from_verilog of Asconp_HPC2_ClockGating_d1 is
  signal SboxInst_n193 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1250
  signal SboxInst_n194 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1249
  signal SboxInst_n195 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1248
  signal SboxInst_n196 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1247
  signal SboxInst_n197 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1246
  signal SboxInst_n198 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1245
  signal SboxInst_n199 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1244
  signal SboxInst_n200 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1243
  signal SboxInst_n201 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1242
  signal SboxInst_n202 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1241
  signal SboxInst_n203 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1240
  signal SboxInst_n204 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1239
  signal SboxInst_n205 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1238
  signal SboxInst_n206 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1237
  signal SboxInst_n207 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1236
  signal SboxInst_n208 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1235
  signal SboxInst_n209 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1234
  signal SboxInst_n210 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1233
  signal SboxInst_n211 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1232
  signal SboxInst_n212 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1231
  signal SboxInst_n213 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1230
  signal SboxInst_n214 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1229
  signal SboxInst_n215 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1228
  signal SboxInst_n216 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1227
  signal SboxInst_n217 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1226
  signal SboxInst_n218 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1225
  signal SboxInst_n219 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1224
  signal SboxInst_n220 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1223
  signal SboxInst_n221 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1222
  signal SboxInst_n222 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1221
  signal SboxInst_n223 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1220
  signal SboxInst_n224 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1219
  signal SboxInst_n225 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1218
  signal SboxInst_n226 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1217
  signal SboxInst_n227 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1216
  signal SboxInst_n228 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1215
  signal SboxInst_n229 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1214
  signal SboxInst_n230 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1213
  signal SboxInst_n231 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1212
  signal SboxInst_n232 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1211
  signal SboxInst_n233 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1210
  signal SboxInst_n234 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1209
  signal SboxInst_n235 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1208
  signal SboxInst_n236 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1207
  signal SboxInst_n237 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1206
  signal SboxInst_n238 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1205
  signal SboxInst_n239 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1204
  signal SboxInst_n240 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1203
  signal SboxInst_n241 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1202
  signal SboxInst_n242 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1201
  signal SboxInst_n243 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1200
  signal SboxInst_n244 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1199
  signal SboxInst_n245 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1198
  signal SboxInst_n246 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1197
  signal SboxInst_n247 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1196
  signal SboxInst_n248 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1195
  signal SboxInst_n249 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1194
  signal SboxInst_n250 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1193
  signal SboxInst_n251 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1192
  signal SboxInst_n252 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1191
  signal SboxInst_n253 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1190
  signal SboxInst_n254 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1189
  signal SboxInst_n255 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1188
  signal SboxInst_n256 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1187
  signal SboxInst_n257 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1186
  signal SboxInst_n258 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1185
  signal SboxInst_n259 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1184
  signal SboxInst_n260 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1183
  signal SboxInst_n261 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1182
  signal SboxInst_n262 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1181
  signal SboxInst_n263 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1180
  signal SboxInst_n264 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1179
  signal SboxInst_n265 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1178
  signal SboxInst_n266 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1177
  signal SboxInst_n267 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1176
  signal SboxInst_n268 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1175
  signal SboxInst_n269 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1174
  signal SboxInst_n270 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1173
  signal SboxInst_n271 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1172
  signal SboxInst_n272 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1171
  signal SboxInst_n273 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1170
  signal SboxInst_n274 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1169
  signal SboxInst_n275 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1168
  signal SboxInst_n276 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1167
  signal SboxInst_n277 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1166
  signal SboxInst_n278 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1165
  signal SboxInst_n279 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1164
  signal SboxInst_n280 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1163
  signal SboxInst_n281 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1162
  signal SboxInst_n282 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1161
  signal SboxInst_n283 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1160
  signal SboxInst_n284 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1159
  signal SboxInst_n285 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1158
  signal SboxInst_n286 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1157
  signal SboxInst_n287 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1156
  signal SboxInst_n288 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1155
  signal SboxInst_n289 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1154
  signal SboxInst_n290 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1153
  signal SboxInst_n291 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1152
  signal SboxInst_n292 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1151
  signal SboxInst_n293 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1150
  signal SboxInst_n294 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1149
  signal SboxInst_n295 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1148
  signal SboxInst_n296 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1147
  signal SboxInst_n297 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1146
  signal SboxInst_n298 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1145
  signal SboxInst_n299 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1144
  signal SboxInst_n300 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1143
  signal SboxInst_n301 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1142
  signal SboxInst_n302 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1141
  signal SboxInst_n303 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1140
  signal SboxInst_n304 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1139
  signal SboxInst_n305 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1138
  signal SboxInst_n306 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1137
  signal SboxInst_n307 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1136
  signal SboxInst_n308 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1135
  signal SboxInst_n309 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1134
  signal SboxInst_n310 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1133
  signal SboxInst_n311 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1132
  signal SboxInst_n312 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1131
  signal SboxInst_n313 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1130
  signal SboxInst_n314 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1129
  signal SboxInst_n315 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1128
  signal SboxInst_n316 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1127
  signal SboxInst_n317 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1126
  signal SboxInst_n318 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1125
  signal SboxInst_n319 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1124
  signal SboxInst_n320 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1123
  signal SboxInst_n321 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1122
  signal SboxInst_n322 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1121
  signal SboxInst_n323 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1120
  signal SboxInst_n324 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1119
  signal SboxInst_n325 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1118
  signal SboxInst_n326 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1117
  signal SboxInst_n327 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1116
  signal SboxInst_n328 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1115
  signal SboxInst_n329 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1114
  signal SboxInst_n330 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1113
  signal SboxInst_n331 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1112
  signal SboxInst_n332 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1111
  signal SboxInst_n333 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1110
  signal SboxInst_n334 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1109
  signal SboxInst_n335 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1108
  signal SboxInst_n336 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1107
  signal SboxInst_n337 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1106
  signal SboxInst_n338 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1105
  signal SboxInst_n339 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1104
  signal SboxInst_n340 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1103
  signal SboxInst_n341 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1102
  signal SboxInst_n342 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1101
  signal SboxInst_n343 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1100
  signal SboxInst_n344 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1099
  signal SboxInst_n345 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1098
  signal SboxInst_n346 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1097
  signal SboxInst_n347 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1096
  signal SboxInst_n348 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1095
  signal SboxInst_n349 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1094
  signal SboxInst_n350 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1093
  signal SboxInst_n351 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1092
  signal SboxInst_n352 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1091
  signal SboxInst_n353 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1090
  signal SboxInst_n354 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1089
  signal SboxInst_n355 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1088
  signal SboxInst_n356 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1087
  signal SboxInst_n357 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1086
  signal SboxInst_n358 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1085
  signal SboxInst_n359 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1084
  signal SboxInst_n360 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1083
  signal SboxInst_n361 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1082
  signal SboxInst_n362 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1081
  signal SboxInst_n363 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1080
  signal SboxInst_n364 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1079
  signal SboxInst_n365 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1078
  signal SboxInst_n366 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1077
  signal SboxInst_n367 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1076
  signal SboxInst_n368 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1075
  signal SboxInst_n369 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1074
  signal SboxInst_n370 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1073
  signal SboxInst_n371 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1072
  signal SboxInst_n372 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1071
  signal SboxInst_n373 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1070
  signal SboxInst_n374 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1069
  signal SboxInst_n375 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1068
  signal SboxInst_n376 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1067
  signal SboxInst_n377 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1066
  signal SboxInst_n378 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1065
  signal SboxInst_n379 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1064
  signal SboxInst_n380 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1063
  signal SboxInst_n381 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1062
  signal SboxInst_n382 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1061
  signal SboxInst_n383 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1060
  signal SboxInst_n384 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1059
  signal tmp_ivl_1 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2940
  signal tmp_ivl_1000 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2974
  signal tmp_ivl_10004 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3461
  signal tmp_ivl_10007 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3461
  signal tmp_ivl_10008 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3461
  signal tmp_ivl_1001 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2974
  signal tmp_ivl_10013 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3461
  signal tmp_ivl_10015 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3461
  signal tmp_ivl_10021 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3462
  signal tmp_ivl_10023 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3462
  signal tmp_ivl_10024 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3462
  signal tmp_ivl_10029 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3462
  signal tmp_ivl_10031 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3462
  signal tmp_ivl_10036 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3462
  signal tmp_ivl_10038 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3462
  signal tmp_ivl_10043 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3463
  signal tmp_ivl_10048 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3463
  signal tmp_ivl_10050 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3463
  signal tmp_ivl_10055 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3463
  signal tmp_ivl_10057 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3463
  signal tmp_ivl_1006 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2974
  signal tmp_ivl_10063 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3464
  signal tmp_ivl_10065 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3464
  signal tmp_ivl_10066 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3464
  signal tmp_ivl_10071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3464
  signal tmp_ivl_10074 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3464
  signal tmp_ivl_10075 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3464
  signal tmp_ivl_1008 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2974
  signal tmp_ivl_10080 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3464
  signal tmp_ivl_10082 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3464
  signal tmp_ivl_10088 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3465
  signal tmp_ivl_10090 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3465
  signal tmp_ivl_10091 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3465
  signal tmp_ivl_10096 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3465
  signal tmp_ivl_10098 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3465
  signal tmp_ivl_101 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2943
  signal tmp_ivl_1010 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2974
  signal tmp_ivl_10103 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3465
  signal tmp_ivl_10105 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3465
  signal tmp_ivl_10110 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3466
  signal tmp_ivl_10115 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3466
  signal tmp_ivl_10117 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3466
  signal tmp_ivl_10122 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3466
  signal tmp_ivl_10124 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3466
  signal tmp_ivl_10126 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3466
  signal tmp_ivl_10128 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3466
  signal tmp_ivl_10134 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3467
  signal tmp_ivl_10135 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3467
  signal tmp_ivl_10140 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3467
  signal tmp_ivl_10143 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3467
  signal tmp_ivl_10145 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3467
  signal tmp_ivl_10146 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3467
  signal tmp_ivl_10151 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3467
  signal tmp_ivl_10153 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3467
  signal tmp_ivl_10159 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3468
  signal tmp_ivl_1016 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2975
  signal tmp_ivl_10160 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3468
  signal tmp_ivl_10165 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3468
  signal tmp_ivl_10167 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3468
  signal tmp_ivl_10172 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3468
  signal tmp_ivl_10174 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3468
  signal tmp_ivl_10179 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3469
  signal tmp_ivl_1018 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2975
  signal tmp_ivl_10184 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3469
  signal tmp_ivl_10186 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3469
  signal tmp_ivl_1019 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2975
  signal tmp_ivl_10191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3469
  signal tmp_ivl_10193 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3469
  signal tmp_ivl_10199 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3470
  signal tmp_ivl_102 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2943
  signal tmp_ivl_10200 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3470
  signal tmp_ivl_10205 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3470
  signal tmp_ivl_10208 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3470
  signal tmp_ivl_10210 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3470
  signal tmp_ivl_10211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3470
  signal tmp_ivl_10216 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3470
  signal tmp_ivl_10218 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3470
  signal tmp_ivl_10224 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3471
  signal tmp_ivl_10225 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3471
  signal tmp_ivl_10230 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3471
  signal tmp_ivl_10233 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3471
  signal tmp_ivl_10235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3471
  signal tmp_ivl_10236 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3471
  signal tmp_ivl_1024 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2975
  signal tmp_ivl_10241 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3471
  signal tmp_ivl_10243 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3471
  signal tmp_ivl_10249 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3472
  signal tmp_ivl_10251 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3472
  signal tmp_ivl_10252 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3472
  signal tmp_ivl_10257 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3472
  signal tmp_ivl_10259 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3472
  signal tmp_ivl_10264 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3472
  signal tmp_ivl_10266 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3472
  signal tmp_ivl_1027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2975
  signal tmp_ivl_10271 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3473
  signal tmp_ivl_10276 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3473
  signal tmp_ivl_10278 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3473
  signal tmp_ivl_10283 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3473
  signal tmp_ivl_10285 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3473
  signal tmp_ivl_1029 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2975
  signal tmp_ivl_10290 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3474
  signal tmp_ivl_10295 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3474
  signal tmp_ivl_10297 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3474
  signal tmp_ivl_1030 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2975
  signal tmp_ivl_10302 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3474
  signal tmp_ivl_10304 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3474
  signal tmp_ivl_10310 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3475
  signal tmp_ivl_10311 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3475
  signal tmp_ivl_10316 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3475
  signal tmp_ivl_10319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3475
  signal tmp_ivl_10321 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3475
  signal tmp_ivl_10322 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3475
  signal tmp_ivl_10327 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3475
  signal tmp_ivl_10329 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3475
  signal tmp_ivl_10335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3476
  signal tmp_ivl_10336 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3476
  signal tmp_ivl_10341 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3476
  signal tmp_ivl_10344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3476
  signal tmp_ivl_10346 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3476
  signal tmp_ivl_10347 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3476
  signal tmp_ivl_1035 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2975
  signal tmp_ivl_10352 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3476
  signal tmp_ivl_10354 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3476
  signal tmp_ivl_10360 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3477
  signal tmp_ivl_10362 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3477
  signal tmp_ivl_10363 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3477
  signal tmp_ivl_10368 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3477
  signal tmp_ivl_1037 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2975
  signal tmp_ivl_10370 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3477
  signal tmp_ivl_10375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3477
  signal tmp_ivl_10377 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3477
  signal tmp_ivl_10382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3478
  signal tmp_ivl_10387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3478
  signal tmp_ivl_10389 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3478
  signal tmp_ivl_1039 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2975
  signal tmp_ivl_10394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3478
  signal tmp_ivl_10396 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3478
  signal tmp_ivl_10401 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3479
  signal tmp_ivl_10406 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3479
  signal tmp_ivl_10408 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3479
  signal tmp_ivl_10413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3479
  signal tmp_ivl_10415 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3479
  signal tmp_ivl_10417 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3479
  signal tmp_ivl_10419 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3479
  signal tmp_ivl_10425 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3480
  signal tmp_ivl_10426 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3480
  signal tmp_ivl_10431 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3480
  signal tmp_ivl_10434 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3480
  signal tmp_ivl_10436 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3480
  signal tmp_ivl_10437 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3480
  signal tmp_ivl_10442 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3480
  signal tmp_ivl_10444 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3480
  signal tmp_ivl_1045 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2976
  signal tmp_ivl_10450 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3481
  signal tmp_ivl_10451 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3481
  signal tmp_ivl_10456 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3481
  signal tmp_ivl_10458 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3481
  signal tmp_ivl_10463 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3481
  signal tmp_ivl_10465 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3481
  signal tmp_ivl_1047 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2976
  signal tmp_ivl_10470 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3482
  signal tmp_ivl_10475 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3482
  signal tmp_ivl_10477 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3482
  signal tmp_ivl_1048 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2976
  signal tmp_ivl_10482 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3482
  signal tmp_ivl_10484 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3482
  signal tmp_ivl_10490 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3483
  signal tmp_ivl_10491 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3483
  signal tmp_ivl_10496 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3483
  signal tmp_ivl_10499 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3483
  signal tmp_ivl_10501 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3483
  signal tmp_ivl_10502 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3483
  signal tmp_ivl_10507 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3483
  signal tmp_ivl_10509 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3483
  signal tmp_ivl_10515 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3484
  signal tmp_ivl_10516 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3484
  signal tmp_ivl_10521 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3484
  signal tmp_ivl_10524 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3484
  signal tmp_ivl_10526 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3484
  signal tmp_ivl_10527 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3484
  signal tmp_ivl_1053 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2976
  signal tmp_ivl_10532 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3484
  signal tmp_ivl_10534 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3484
  signal tmp_ivl_10540 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3485
  signal tmp_ivl_10542 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3485
  signal tmp_ivl_10543 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3485
  signal tmp_ivl_10548 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3485
  signal tmp_ivl_10550 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3485
  signal tmp_ivl_10555 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3485
  signal tmp_ivl_10557 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3485
  signal tmp_ivl_1056 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2976
  signal tmp_ivl_10562 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3486
  signal tmp_ivl_10567 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3486
  signal tmp_ivl_10569 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3486
  signal tmp_ivl_10574 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3486
  signal tmp_ivl_10576 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3486
  signal tmp_ivl_1058 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2976
  signal tmp_ivl_10581 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3487
  signal tmp_ivl_10586 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3487
  signal tmp_ivl_10588 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3487
  signal tmp_ivl_1059 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2976
  signal tmp_ivl_10593 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3487
  signal tmp_ivl_10595 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3487
  signal tmp_ivl_10601 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3488
  signal tmp_ivl_10602 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3488
  signal tmp_ivl_10607 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3488
  signal tmp_ivl_10610 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3488
  signal tmp_ivl_10612 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3488
  signal tmp_ivl_10613 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3488
  signal tmp_ivl_10618 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3488
  signal tmp_ivl_10620 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3488
  signal tmp_ivl_10626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3489
  signal tmp_ivl_10627 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3489
  signal tmp_ivl_10632 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3489
  signal tmp_ivl_10635 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3489
  signal tmp_ivl_10637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3489
  signal tmp_ivl_10638 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3489
  signal tmp_ivl_1064 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2976
  signal tmp_ivl_10643 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3489
  signal tmp_ivl_10645 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3489
  signal tmp_ivl_10651 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3490
  signal tmp_ivl_10653 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3490
  signal tmp_ivl_10654 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3490
  signal tmp_ivl_10659 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3490
  signal tmp_ivl_1066 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2976
  signal tmp_ivl_10661 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3490
  signal tmp_ivl_10666 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3490
  signal tmp_ivl_10668 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3490
  signal tmp_ivl_10673 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3491
  signal tmp_ivl_10678 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3491
  signal tmp_ivl_1068 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2976
  signal tmp_ivl_10680 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3491
  signal tmp_ivl_10685 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3491
  signal tmp_ivl_10687 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3491
  signal tmp_ivl_10692 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3492
  signal tmp_ivl_10697 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3492
  signal tmp_ivl_10699 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3492
  signal tmp_ivl_107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2943
  signal tmp_ivl_10704 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3492
  signal tmp_ivl_10706 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3492
  signal tmp_ivl_10708 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3492
  signal tmp_ivl_10710 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3492
  signal tmp_ivl_10715 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3493
  signal tmp_ivl_10720 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3493
  signal tmp_ivl_10722 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3493
  signal tmp_ivl_10727 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3493
  signal tmp_ivl_10729 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3493
  signal tmp_ivl_10735 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3494
  signal tmp_ivl_10737 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3494
  signal tmp_ivl_10738 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3494
  signal tmp_ivl_1074 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2977
  signal tmp_ivl_10743 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3494
  signal tmp_ivl_10746 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3494
  signal tmp_ivl_10747 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3494
  signal tmp_ivl_10752 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3494
  signal tmp_ivl_10754 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3494
  signal tmp_ivl_1076 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2977
  signal tmp_ivl_10760 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3495
  signal tmp_ivl_10762 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3495
  signal tmp_ivl_10763 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3495
  signal tmp_ivl_10768 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3495
  signal tmp_ivl_1077 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2977
  signal tmp_ivl_10770 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3495
  signal tmp_ivl_10775 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3495
  signal tmp_ivl_10777 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3495
  signal tmp_ivl_10782 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3496
  signal tmp_ivl_10787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3496
  signal tmp_ivl_10789 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3496
  signal tmp_ivl_10794 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3496
  signal tmp_ivl_10796 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3496
  signal tmp_ivl_10798 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3496
  signal tmp_ivl_10800 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3496
  signal tmp_ivl_10805 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3497
  signal tmp_ivl_10810 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3497
  signal tmp_ivl_10812 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3497
  signal tmp_ivl_10817 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3497
  signal tmp_ivl_10819 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3497
  signal tmp_ivl_1082 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2977
  signal tmp_ivl_10825 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3498
  signal tmp_ivl_10827 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3498
  signal tmp_ivl_10828 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3498
  signal tmp_ivl_10833 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3498
  signal tmp_ivl_10836 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3498
  signal tmp_ivl_10837 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3498
  signal tmp_ivl_10842 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3498
  signal tmp_ivl_10844 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3498
  signal tmp_ivl_1085 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2977
  signal tmp_ivl_10850 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3499
  signal tmp_ivl_10852 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3499
  signal tmp_ivl_10853 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3499
  signal tmp_ivl_10858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3499
  signal tmp_ivl_10860 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3499
  signal tmp_ivl_10865 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3499
  signal tmp_ivl_10867 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3499
  signal tmp_ivl_1087 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2977
  signal tmp_ivl_10872 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3500
  signal tmp_ivl_10877 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3500
  signal tmp_ivl_10879 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3500
  signal tmp_ivl_1088 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2977
  signal tmp_ivl_10884 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3500
  signal tmp_ivl_10886 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3500
  signal tmp_ivl_10888 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3500
  signal tmp_ivl_10890 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3500
  signal tmp_ivl_10896 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3501
  signal tmp_ivl_10898 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3501
  signal tmp_ivl_10899 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3501
  signal tmp_ivl_109 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2943
  signal tmp_ivl_10904 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3501
  signal tmp_ivl_10907 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3501
  signal tmp_ivl_10908 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3501
  signal tmp_ivl_10913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3501
  signal tmp_ivl_10915 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3501
  signal tmp_ivl_10921 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3502
  signal tmp_ivl_10923 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3502
  signal tmp_ivl_10924 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3502
  signal tmp_ivl_10929 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3502
  signal tmp_ivl_1093 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2977
  signal tmp_ivl_10931 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3502
  signal tmp_ivl_10936 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3502
  signal tmp_ivl_10938 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3502
  signal tmp_ivl_10943 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3503
  signal tmp_ivl_10948 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3503
  signal tmp_ivl_1095 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2977
  signal tmp_ivl_10950 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3503
  signal tmp_ivl_10955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3503
  signal tmp_ivl_10957 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3503
  signal tmp_ivl_10963 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3504
  signal tmp_ivl_10965 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3504
  signal tmp_ivl_10966 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3504
  signal tmp_ivl_1097 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2977
  signal tmp_ivl_10971 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3504
  signal tmp_ivl_10974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3504
  signal tmp_ivl_10975 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3504
  signal tmp_ivl_10980 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3504
  signal tmp_ivl_10982 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3504
  signal tmp_ivl_10988 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3505
  signal tmp_ivl_10990 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3505
  signal tmp_ivl_10991 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3505
  signal tmp_ivl_10996 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3505
  signal tmp_ivl_10998 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3505
  signal tmp_ivl_11003 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3505
  signal tmp_ivl_11005 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3505
  signal tmp_ivl_11010 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3506
  signal tmp_ivl_11015 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3506
  signal tmp_ivl_11017 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3506
  signal tmp_ivl_11022 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3506
  signal tmp_ivl_11024 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3506
  signal tmp_ivl_11026 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3506
  signal tmp_ivl_11028 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3506
  signal tmp_ivl_1103 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2978
  signal tmp_ivl_11034 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3507
  signal tmp_ivl_11035 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3507
  signal tmp_ivl_11040 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3507
  signal tmp_ivl_11043 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3507
  signal tmp_ivl_11045 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3507
  signal tmp_ivl_11046 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3507
  signal tmp_ivl_1105 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2978
  signal tmp_ivl_11051 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3507
  signal tmp_ivl_11053 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3507
  signal tmp_ivl_11059 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3508
  signal tmp_ivl_1106 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2978
  signal tmp_ivl_11060 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3508
  signal tmp_ivl_11065 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3508
  signal tmp_ivl_11068 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3508
  signal tmp_ivl_11070 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3508
  signal tmp_ivl_11071 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3508
  signal tmp_ivl_11076 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3508
  signal tmp_ivl_11078 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3508
  signal tmp_ivl_11084 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3509
  signal tmp_ivl_11086 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3509
  signal tmp_ivl_11087 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3509
  signal tmp_ivl_11092 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3509
  signal tmp_ivl_11094 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3509
  signal tmp_ivl_11099 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3509
  signal tmp_ivl_111 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2943
  signal tmp_ivl_11101 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3509
  signal tmp_ivl_11106 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3510
  signal tmp_ivl_1111 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2978
  signal tmp_ivl_11111 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3510
  signal tmp_ivl_11113 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3510
  signal tmp_ivl_11118 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3510
  signal tmp_ivl_11120 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3510
  signal tmp_ivl_11126 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3511
  signal tmp_ivl_11127 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3511
  signal tmp_ivl_11132 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3511
  signal tmp_ivl_11135 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3511
  signal tmp_ivl_11137 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3511
  signal tmp_ivl_11138 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3511
  signal tmp_ivl_1114 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2978
  signal tmp_ivl_11143 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3511
  signal tmp_ivl_11145 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3511
  signal tmp_ivl_11151 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3512
  signal tmp_ivl_11152 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3512
  signal tmp_ivl_11157 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3512
  signal tmp_ivl_11159 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3512
  signal tmp_ivl_1116 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2978
  signal tmp_ivl_11164 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3512
  signal tmp_ivl_11166 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3512
  signal tmp_ivl_1117 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2978
  signal tmp_ivl_11171 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3513
  signal tmp_ivl_11176 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3513
  signal tmp_ivl_11178 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3513
  signal tmp_ivl_11183 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3513
  signal tmp_ivl_11185 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3513
  signal tmp_ivl_11190 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3514
  signal tmp_ivl_11195 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3514
  signal tmp_ivl_11197 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3514
  signal tmp_ivl_11202 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3514
  signal tmp_ivl_11204 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3514
  signal tmp_ivl_11210 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3515
  signal tmp_ivl_11211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3515
  signal tmp_ivl_11216 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3515
  signal tmp_ivl_11219 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3515
  signal tmp_ivl_1122 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2978
  signal tmp_ivl_11221 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3515
  signal tmp_ivl_11222 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3515
  signal tmp_ivl_11227 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3515
  signal tmp_ivl_11229 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3515
  signal tmp_ivl_11235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3516
  signal tmp_ivl_11236 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3516
  signal tmp_ivl_1124 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2978
  signal tmp_ivl_11241 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3516
  signal tmp_ivl_11244 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3516
  signal tmp_ivl_11246 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3516
  signal tmp_ivl_11247 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3516
  signal tmp_ivl_11252 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3516
  signal tmp_ivl_11254 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3516
  signal tmp_ivl_1126 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2978
  signal tmp_ivl_11260 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3517
  signal tmp_ivl_11262 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3517
  signal tmp_ivl_11263 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3517
  signal tmp_ivl_11268 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3517
  signal tmp_ivl_11270 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3517
  signal tmp_ivl_11275 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3517
  signal tmp_ivl_11277 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3517
  signal tmp_ivl_11282 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3518
  signal tmp_ivl_11287 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3518
  signal tmp_ivl_11289 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3518
  signal tmp_ivl_11294 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3518
  signal tmp_ivl_11296 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3518
  signal tmp_ivl_11301 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3519
  signal tmp_ivl_11306 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3519
  signal tmp_ivl_11308 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3519
  signal tmp_ivl_11313 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3519
  signal tmp_ivl_11315 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3519
  signal tmp_ivl_11317 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3519
  signal tmp_ivl_11319 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3519
  signal tmp_ivl_1132 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2979
  signal tmp_ivl_11325 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3520
  signal tmp_ivl_11326 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3520
  signal tmp_ivl_11331 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3520
  signal tmp_ivl_11334 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3520
  signal tmp_ivl_11336 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3520
  signal tmp_ivl_11337 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3520
  signal tmp_ivl_1134 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2979
  signal tmp_ivl_11342 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3520
  signal tmp_ivl_11344 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3520
  signal tmp_ivl_1135 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2979
  signal tmp_ivl_11350 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3521
  signal tmp_ivl_11351 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3521
  signal tmp_ivl_11356 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3521
  signal tmp_ivl_11359 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3521
  signal tmp_ivl_11361 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3521
  signal tmp_ivl_11362 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3521
  signal tmp_ivl_11367 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3521
  signal tmp_ivl_11369 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3521
  signal tmp_ivl_11375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3522
  signal tmp_ivl_11377 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3522
  signal tmp_ivl_11378 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3522
  signal tmp_ivl_11383 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3522
  signal tmp_ivl_11385 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3522
  signal tmp_ivl_11390 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3522
  signal tmp_ivl_11392 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3522
  signal tmp_ivl_11397 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3523
  signal tmp_ivl_1140 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2979
  signal tmp_ivl_11402 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3523
  signal tmp_ivl_11404 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3523
  signal tmp_ivl_11409 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3523
  signal tmp_ivl_11411 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3523
  signal tmp_ivl_11416 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3524
  signal tmp_ivl_11421 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3524
  signal tmp_ivl_11423 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3524
  signal tmp_ivl_11428 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3524
  signal tmp_ivl_1143 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2979
  signal tmp_ivl_11430 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3524
  signal tmp_ivl_11436 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3525
  signal tmp_ivl_11437 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3525
  signal tmp_ivl_11442 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3525
  signal tmp_ivl_11445 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3525
  signal tmp_ivl_11447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3525
  signal tmp_ivl_11448 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3525
  signal tmp_ivl_1145 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2979
  signal tmp_ivl_11453 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3525
  signal tmp_ivl_11455 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3525
  signal tmp_ivl_1146 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2979
  signal tmp_ivl_11461 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3526
  signal tmp_ivl_11462 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3526
  signal tmp_ivl_11467 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3526
  signal tmp_ivl_11469 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3526
  signal tmp_ivl_11474 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3526
  signal tmp_ivl_11476 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3526
  signal tmp_ivl_11481 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3527
  signal tmp_ivl_11486 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3527
  signal tmp_ivl_11488 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3527
  signal tmp_ivl_11493 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3527
  signal tmp_ivl_11495 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3527
  signal tmp_ivl_11500 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3528
  signal tmp_ivl_11505 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3528
  signal tmp_ivl_11507 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3528
  signal tmp_ivl_1151 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2979
  signal tmp_ivl_11512 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3528
  signal tmp_ivl_11514 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3528
  signal tmp_ivl_11516 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3528
  signal tmp_ivl_11518 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3528
  signal tmp_ivl_11524 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3529
  signal tmp_ivl_11525 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3529
  signal tmp_ivl_1153 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2979
  signal tmp_ivl_11530 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3529
  signal tmp_ivl_11533 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3529
  signal tmp_ivl_11535 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3529
  signal tmp_ivl_11536 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3529
  signal tmp_ivl_11541 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3529
  signal tmp_ivl_11543 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3529
  signal tmp_ivl_11549 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3530
  signal tmp_ivl_1155 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2979
  signal tmp_ivl_11550 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3530
  signal tmp_ivl_11555 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3530
  signal tmp_ivl_11558 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3530
  signal tmp_ivl_11560 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3530
  signal tmp_ivl_11561 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3530
  signal tmp_ivl_11566 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3530
  signal tmp_ivl_11568 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3530
  signal tmp_ivl_11574 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3531
  signal tmp_ivl_11576 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3531
  signal tmp_ivl_11577 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3531
  signal tmp_ivl_11582 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3531
  signal tmp_ivl_11584 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3531
  signal tmp_ivl_11589 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3531
  signal tmp_ivl_11591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3531
  signal tmp_ivl_11596 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3532
  signal tmp_ivl_11601 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3532
  signal tmp_ivl_11603 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3532
  signal tmp_ivl_11608 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3532
  signal tmp_ivl_1161 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2980
  signal tmp_ivl_11610 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3532
  signal tmp_ivl_11615 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3533
  signal tmp_ivl_11620 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3533
  signal tmp_ivl_11622 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3533
  signal tmp_ivl_11627 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3533
  signal tmp_ivl_11629 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3533
  signal tmp_ivl_1163 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2980
  signal tmp_ivl_11635 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3534
  signal tmp_ivl_11636 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3534
  signal tmp_ivl_1164 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2980
  signal tmp_ivl_11641 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3534
  signal tmp_ivl_11644 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3534
  signal tmp_ivl_11646 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3534
  signal tmp_ivl_11647 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3534
  signal tmp_ivl_11652 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3534
  signal tmp_ivl_11654 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3534
  signal tmp_ivl_11660 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3535
  signal tmp_ivl_11661 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3535
  signal tmp_ivl_11666 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3535
  signal tmp_ivl_11669 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3535
  signal tmp_ivl_11671 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3535
  signal tmp_ivl_11672 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3535
  signal tmp_ivl_11677 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3535
  signal tmp_ivl_11679 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3535
  signal tmp_ivl_11685 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3536
  signal tmp_ivl_11687 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3536
  signal tmp_ivl_11688 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3536
  signal tmp_ivl_1169 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2980
  signal tmp_ivl_11693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3536
  signal tmp_ivl_11695 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3536
  signal tmp_ivl_117 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2944
  signal tmp_ivl_11700 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3536
  signal tmp_ivl_11702 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3536
  signal tmp_ivl_11707 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3537
  signal tmp_ivl_11712 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3537
  signal tmp_ivl_11714 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3537
  signal tmp_ivl_11719 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3537
  signal tmp_ivl_1172 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2980
  signal tmp_ivl_11721 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3537
  signal tmp_ivl_11726 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3538
  signal tmp_ivl_11731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3538
  signal tmp_ivl_11733 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3538
  signal tmp_ivl_11738 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3538
  signal tmp_ivl_1174 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2980
  signal tmp_ivl_11740 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3538
  signal tmp_ivl_11742 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3538
  signal tmp_ivl_11744 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3538
  signal tmp_ivl_11749 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3539
  signal tmp_ivl_1175 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2980
  signal tmp_ivl_11754 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3539
  signal tmp_ivl_11756 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3539
  signal tmp_ivl_11761 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3539
  signal tmp_ivl_11763 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3539
  signal tmp_ivl_11769 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3540
  signal tmp_ivl_11771 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3540
  signal tmp_ivl_11772 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3540
  signal tmp_ivl_11777 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3540
  signal tmp_ivl_11780 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3540
  signal tmp_ivl_11781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3540
  signal tmp_ivl_11786 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3540
  signal tmp_ivl_11788 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3540
  signal tmp_ivl_11794 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3541
  signal tmp_ivl_11796 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3541
  signal tmp_ivl_11797 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3541
  signal tmp_ivl_1180 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2980
  signal tmp_ivl_11802 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3541
  signal tmp_ivl_11804 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3541
  signal tmp_ivl_11809 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3541
  signal tmp_ivl_11811 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3541
  signal tmp_ivl_11816 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3542
  signal tmp_ivl_1182 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2980
  signal tmp_ivl_11821 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3542
  signal tmp_ivl_11823 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3542
  signal tmp_ivl_11828 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3542
  signal tmp_ivl_11830 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3542
  signal tmp_ivl_11832 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3542
  signal tmp_ivl_11834 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3542
  signal tmp_ivl_11839 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3543
  signal tmp_ivl_1184 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2980
  signal tmp_ivl_11844 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3543
  signal tmp_ivl_11846 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3543
  signal tmp_ivl_11851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3543
  signal tmp_ivl_11853 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3543
  signal tmp_ivl_11858 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3544
  signal tmp_ivl_11863 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3544
  signal tmp_ivl_11865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3544
  signal tmp_ivl_11870 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3544
  signal tmp_ivl_11872 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3544
  signal tmp_ivl_11874 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3544
  signal tmp_ivl_11876 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3544
  signal tmp_ivl_11882 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3545
  signal tmp_ivl_11883 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3545
  signal tmp_ivl_11888 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3545
  signal tmp_ivl_11891 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3545
  signal tmp_ivl_11893 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3545
  signal tmp_ivl_11894 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3545
  signal tmp_ivl_11899 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3545
  signal tmp_ivl_119 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2944
  signal tmp_ivl_1190 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2981
  signal tmp_ivl_11901 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3545
  signal tmp_ivl_11907 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3546
  signal tmp_ivl_11908 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3546
  signal tmp_ivl_11913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3546
  signal tmp_ivl_11916 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3546
  signal tmp_ivl_11918 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3546
  signal tmp_ivl_11919 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3546
  signal tmp_ivl_1192 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2981
  signal tmp_ivl_11924 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3546
  signal tmp_ivl_11926 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3546
  signal tmp_ivl_1193 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2981
  signal tmp_ivl_11932 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3547
  signal tmp_ivl_11934 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3547
  signal tmp_ivl_11935 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3547
  signal tmp_ivl_11940 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3547
  signal tmp_ivl_11942 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3547
  signal tmp_ivl_11947 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3547
  signal tmp_ivl_11949 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3547
  signal tmp_ivl_11954 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3548
  signal tmp_ivl_11959 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3548
  signal tmp_ivl_11961 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3548
  signal tmp_ivl_11966 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3548
  signal tmp_ivl_11968 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3548
  signal tmp_ivl_11973 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3549
  signal tmp_ivl_11978 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3549
  signal tmp_ivl_1198 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2981
  signal tmp_ivl_11980 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3549
  signal tmp_ivl_11985 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3549
  signal tmp_ivl_11987 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3549
  signal tmp_ivl_11993 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3550
  signal tmp_ivl_11994 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3550
  signal tmp_ivl_11999 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3550
  signal tmp_ivl_12 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2940
  signal tmp_ivl_120 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2944
  signal tmp_ivl_12002 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3550
  signal tmp_ivl_12004 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3550
  signal tmp_ivl_12005 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3550
  signal tmp_ivl_1201 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2981
  signal tmp_ivl_12010 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3550
  signal tmp_ivl_12012 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3550
  signal tmp_ivl_12018 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3551
  signal tmp_ivl_12019 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3551
  signal tmp_ivl_12024 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3551
  signal tmp_ivl_12026 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3551
  signal tmp_ivl_1203 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2981
  signal tmp_ivl_12031 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3551
  signal tmp_ivl_12033 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3551
  signal tmp_ivl_12038 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3552
  signal tmp_ivl_1204 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2981
  signal tmp_ivl_12043 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3552
  signal tmp_ivl_12045 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3552
  signal tmp_ivl_12050 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3552
  signal tmp_ivl_12052 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3552
  signal tmp_ivl_12057 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3553
  signal tmp_ivl_12062 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3553
  signal tmp_ivl_12064 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3553
  signal tmp_ivl_12069 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3553
  signal tmp_ivl_12071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3553
  signal tmp_ivl_12073 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3553
  signal tmp_ivl_12075 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3553
  signal tmp_ivl_12080 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3554
  signal tmp_ivl_12085 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3554
  signal tmp_ivl_12087 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3554
  signal tmp_ivl_1209 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2981
  signal tmp_ivl_12092 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3554
  signal tmp_ivl_12094 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3554
  signal tmp_ivl_12100 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3555
  signal tmp_ivl_12102 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3555
  signal tmp_ivl_12103 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3555
  signal tmp_ivl_12108 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3555
  signal tmp_ivl_1211 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2981
  signal tmp_ivl_12111 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3555
  signal tmp_ivl_12112 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3555
  signal tmp_ivl_12117 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3555
  signal tmp_ivl_12119 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3555
  signal tmp_ivl_12125 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3556
  signal tmp_ivl_12127 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3556
  signal tmp_ivl_12128 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3556
  signal tmp_ivl_1213 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2981
  signal tmp_ivl_12133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3556
  signal tmp_ivl_12135 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3556
  signal tmp_ivl_12140 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3556
  signal tmp_ivl_12142 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3556
  signal tmp_ivl_12147 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3557
  signal tmp_ivl_12152 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3557
  signal tmp_ivl_12154 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3557
  signal tmp_ivl_12159 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3557
  signal tmp_ivl_12161 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3557
  signal tmp_ivl_12163 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3557
  signal tmp_ivl_12165 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3557
  signal tmp_ivl_12171 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3558
  signal tmp_ivl_12172 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3558
  signal tmp_ivl_12177 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3558
  signal tmp_ivl_12180 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3558
  signal tmp_ivl_12182 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3558
  signal tmp_ivl_12183 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3558
  signal tmp_ivl_12188 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3558
  signal tmp_ivl_1219 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2982
  signal tmp_ivl_12190 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3558
  signal tmp_ivl_12195 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3559
  signal tmp_ivl_12200 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3559
  signal tmp_ivl_12202 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3559
  signal tmp_ivl_12207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3559
  signal tmp_ivl_12209 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3559
  signal tmp_ivl_1221 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2982
  signal tmp_ivl_12215 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3560
  signal tmp_ivl_12216 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3560
  signal tmp_ivl_1222 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2982
  signal tmp_ivl_12221 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3560
  signal tmp_ivl_12224 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3560
  signal tmp_ivl_12226 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3560
  signal tmp_ivl_12227 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3560
  signal tmp_ivl_12232 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3560
  signal tmp_ivl_12234 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3560
  signal tmp_ivl_12239 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3561
  signal tmp_ivl_12244 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3561
  signal tmp_ivl_12246 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3561
  signal tmp_ivl_12251 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3561
  signal tmp_ivl_12253 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3561
  signal tmp_ivl_12258 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3562
  signal tmp_ivl_12263 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3562
  signal tmp_ivl_12265 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3562
  signal tmp_ivl_1227 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2982
  signal tmp_ivl_12270 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3562
  signal tmp_ivl_12272 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3562
  signal tmp_ivl_12277 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3563
  signal tmp_ivl_12282 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3563
  signal tmp_ivl_12284 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3563
  signal tmp_ivl_12289 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3563
  signal tmp_ivl_12291 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3563
  signal tmp_ivl_12296 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3564
  signal tmp_ivl_1230 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2982
  signal tmp_ivl_12301 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3564
  signal tmp_ivl_12303 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3564
  signal tmp_ivl_12308 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3564
  signal tmp_ivl_12310 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3564
  signal tmp_ivl_12312 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3564
  signal tmp_ivl_12314 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3564
  signal tmp_ivl_1232 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2982
  signal tmp_ivl_12320 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3565
  signal tmp_ivl_12322 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3565
  signal tmp_ivl_12323 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3565
  signal tmp_ivl_12328 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3565
  signal tmp_ivl_1233 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2982
  signal tmp_ivl_12331 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3565
  signal tmp_ivl_12332 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3565
  signal tmp_ivl_12337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3565
  signal tmp_ivl_12339 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3565
  signal tmp_ivl_12345 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3566
  signal tmp_ivl_12347 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3566
  signal tmp_ivl_12348 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3566
  signal tmp_ivl_12353 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3566
  signal tmp_ivl_12355 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3566
  signal tmp_ivl_12360 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3566
  signal tmp_ivl_12362 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3566
  signal tmp_ivl_12367 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3567
  signal tmp_ivl_12372 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3567
  signal tmp_ivl_12374 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3567
  signal tmp_ivl_12379 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3567
  signal tmp_ivl_1238 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2982
  signal tmp_ivl_12381 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3567
  signal tmp_ivl_12387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3568
  signal tmp_ivl_12389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3568
  signal tmp_ivl_12390 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3568
  signal tmp_ivl_12395 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3568
  signal tmp_ivl_12398 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3568
  signal tmp_ivl_12399 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3568
  signal tmp_ivl_1240 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2982
  signal tmp_ivl_12404 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3568
  signal tmp_ivl_12406 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3568
  signal tmp_ivl_12412 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3569
  signal tmp_ivl_12414 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3569
  signal tmp_ivl_12415 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3569
  signal tmp_ivl_1242 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2982
  signal tmp_ivl_12420 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3569
  signal tmp_ivl_12422 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3569
  signal tmp_ivl_12427 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3569
  signal tmp_ivl_12429 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3569
  signal tmp_ivl_12434 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3570
  signal tmp_ivl_12439 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3570
  signal tmp_ivl_12441 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3570
  signal tmp_ivl_12446 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3570
  signal tmp_ivl_12448 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3570
  signal tmp_ivl_12450 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3570
  signal tmp_ivl_12452 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3570
  signal tmp_ivl_12457 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3571
  signal tmp_ivl_12462 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3571
  signal tmp_ivl_12464 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3571
  signal tmp_ivl_12469 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3571
  signal tmp_ivl_12471 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3571
  signal tmp_ivl_12476 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3572
  signal tmp_ivl_1248 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2983
  signal tmp_ivl_12481 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3572
  signal tmp_ivl_12483 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3572
  signal tmp_ivl_12488 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3572
  signal tmp_ivl_12490 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3572
  signal tmp_ivl_12492 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3572
  signal tmp_ivl_12494 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3572
  signal tmp_ivl_12499 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3573
  signal tmp_ivl_125 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2944
  signal tmp_ivl_1250 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2983
  signal tmp_ivl_12504 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3573
  signal tmp_ivl_12506 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3573
  signal tmp_ivl_1251 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2983
  signal tmp_ivl_12511 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3573
  signal tmp_ivl_12513 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3573
  signal tmp_ivl_12519 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3574
  signal tmp_ivl_12521 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3574
  signal tmp_ivl_12522 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3574
  signal tmp_ivl_12527 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3574
  signal tmp_ivl_12530 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3574
  signal tmp_ivl_12531 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3574
  signal tmp_ivl_12536 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3574
  signal tmp_ivl_12538 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3574
  signal tmp_ivl_12544 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3575
  signal tmp_ivl_12546 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3575
  signal tmp_ivl_12547 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3575
  signal tmp_ivl_12552 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3575
  signal tmp_ivl_12554 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3575
  signal tmp_ivl_12559 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3575
  signal tmp_ivl_1256 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2983
  signal tmp_ivl_12561 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3575
  signal tmp_ivl_12566 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3576
  signal tmp_ivl_12571 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3576
  signal tmp_ivl_12573 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3576
  signal tmp_ivl_12578 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3576
  signal tmp_ivl_12580 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3576
  signal tmp_ivl_12582 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3576
  signal tmp_ivl_12584 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3576
  signal tmp_ivl_1259 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2983
  signal tmp_ivl_12590 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3577
  signal tmp_ivl_12591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3577
  signal tmp_ivl_12596 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3577
  signal tmp_ivl_12599 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3577
  signal tmp_ivl_12601 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3577
  signal tmp_ivl_12602 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3577
  signal tmp_ivl_12607 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3577
  signal tmp_ivl_12609 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3577
  signal tmp_ivl_1261 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2983
  signal tmp_ivl_12615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3578
  signal tmp_ivl_12616 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3578
  signal tmp_ivl_1262 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2983
  signal tmp_ivl_12621 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3578
  signal tmp_ivl_12624 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3578
  signal tmp_ivl_12626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3578
  signal tmp_ivl_12627 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3578
  signal tmp_ivl_12632 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3578
  signal tmp_ivl_12634 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3578
  signal tmp_ivl_12640 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3579
  signal tmp_ivl_12642 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3579
  signal tmp_ivl_12643 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3579
  signal tmp_ivl_12648 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3579
  signal tmp_ivl_12650 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3579
  signal tmp_ivl_12655 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3579
  signal tmp_ivl_12657 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3579
  signal tmp_ivl_12662 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3580
  signal tmp_ivl_12667 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3580
  signal tmp_ivl_12669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3580
  signal tmp_ivl_1267 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2983
  signal tmp_ivl_12674 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3580
  signal tmp_ivl_12676 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3580
  signal tmp_ivl_12681 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3581
  signal tmp_ivl_12686 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3581
  signal tmp_ivl_12688 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3581
  signal tmp_ivl_1269 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2983
  signal tmp_ivl_12693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3581
  signal tmp_ivl_12695 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3581
  signal tmp_ivl_12701 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3582
  signal tmp_ivl_12702 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3582
  signal tmp_ivl_12707 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3582
  signal tmp_ivl_1271 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2983
  signal tmp_ivl_12710 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3582
  signal tmp_ivl_12712 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3582
  signal tmp_ivl_12713 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3582
  signal tmp_ivl_12718 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3582
  signal tmp_ivl_12720 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3582
  signal tmp_ivl_12726 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3583
  signal tmp_ivl_12727 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3583
  signal tmp_ivl_12732 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3583
  signal tmp_ivl_12735 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3583
  signal tmp_ivl_12737 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3583
  signal tmp_ivl_12738 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3583
  signal tmp_ivl_12743 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3583
  signal tmp_ivl_12745 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3583
  signal tmp_ivl_12751 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3584
  signal tmp_ivl_12753 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3584
  signal tmp_ivl_12754 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3584
  signal tmp_ivl_12759 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3584
  signal tmp_ivl_12761 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3584
  signal tmp_ivl_12766 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3584
  signal tmp_ivl_12768 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3584
  signal tmp_ivl_1277 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2984
  signal tmp_ivl_12773 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3585
  signal tmp_ivl_12778 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3585
  signal tmp_ivl_12780 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3585
  signal tmp_ivl_12785 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3585
  signal tmp_ivl_12787 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3585
  signal tmp_ivl_1279 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2984
  signal tmp_ivl_12792 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3586
  signal tmp_ivl_12797 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3586
  signal tmp_ivl_12799 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3586
  signal tmp_ivl_128 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2944
  signal tmp_ivl_1280 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2984
  signal tmp_ivl_12804 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3586
  signal tmp_ivl_12806 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3586
  signal tmp_ivl_12808 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3586
  signal tmp_ivl_12810 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3586
  signal tmp_ivl_12816 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3587
  signal tmp_ivl_12817 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3587
  signal tmp_ivl_12822 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3587
  signal tmp_ivl_12825 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3587
  signal tmp_ivl_12827 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3587
  signal tmp_ivl_12828 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3587
  signal tmp_ivl_12833 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3587
  signal tmp_ivl_12835 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3587
  signal tmp_ivl_12841 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3588
  signal tmp_ivl_12842 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3588
  signal tmp_ivl_12847 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3588
  signal tmp_ivl_12849 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3588
  signal tmp_ivl_1285 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2984
  signal tmp_ivl_12854 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3588
  signal tmp_ivl_12856 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3588
  signal tmp_ivl_12861 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3589
  signal tmp_ivl_12866 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3589
  signal tmp_ivl_12868 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3589
  signal tmp_ivl_12873 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3589
  signal tmp_ivl_12875 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3589
  signal tmp_ivl_1288 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2984
  signal tmp_ivl_12881 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3590
  signal tmp_ivl_12882 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3590
  signal tmp_ivl_12887 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3590
  signal tmp_ivl_12889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3590
  signal tmp_ivl_12894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3590
  signal tmp_ivl_12896 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3590
  signal tmp_ivl_1290 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2984
  signal tmp_ivl_12901 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3591
  signal tmp_ivl_12906 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3591
  signal tmp_ivl_12908 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3591
  signal tmp_ivl_1291 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2984
  signal tmp_ivl_12913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3591
  signal tmp_ivl_12915 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3591
  signal tmp_ivl_12920 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3592
  signal tmp_ivl_12925 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3592
  signal tmp_ivl_12927 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3592
  signal tmp_ivl_12932 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3592
  signal tmp_ivl_12934 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3592
  signal tmp_ivl_12940 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3593
  signal tmp_ivl_12941 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3593
  signal tmp_ivl_12946 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3593
  signal tmp_ivl_12949 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3593
  signal tmp_ivl_12951 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3593
  signal tmp_ivl_12952 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3593
  signal tmp_ivl_12957 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3593
  signal tmp_ivl_12959 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3593
  signal tmp_ivl_1296 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2984
  signal tmp_ivl_12965 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3594
  signal tmp_ivl_12966 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3594
  signal tmp_ivl_12971 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3594
  signal tmp_ivl_12974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3594
  signal tmp_ivl_12976 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3594
  signal tmp_ivl_12977 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3594
  signal tmp_ivl_1298 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2984
  signal tmp_ivl_12982 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3594
  signal tmp_ivl_12984 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3594
  signal tmp_ivl_12990 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3595
  signal tmp_ivl_12992 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3595
  signal tmp_ivl_12993 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3595
  signal tmp_ivl_12998 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3595
  signal tmp_ivl_130 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2944
  signal tmp_ivl_1300 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2984
  signal tmp_ivl_13000 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3595
  signal tmp_ivl_13005 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3595
  signal tmp_ivl_13007 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3595
  signal tmp_ivl_13012 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3596
  signal tmp_ivl_13017 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3596
  signal tmp_ivl_13019 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3596
  signal tmp_ivl_13024 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3596
  signal tmp_ivl_13026 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3596
  signal tmp_ivl_13031 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3597
  signal tmp_ivl_13036 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3597
  signal tmp_ivl_13038 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3597
  signal tmp_ivl_13043 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3597
  signal tmp_ivl_13045 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3597
  signal tmp_ivl_13047 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3597
  signal tmp_ivl_13049 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3597
  signal tmp_ivl_13054 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3598
  signal tmp_ivl_13059 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3598
  signal tmp_ivl_1306 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2985
  signal tmp_ivl_13061 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3598
  signal tmp_ivl_13066 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3598
  signal tmp_ivl_13068 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3598
  signal tmp_ivl_13074 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3599
  signal tmp_ivl_13076 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3599
  signal tmp_ivl_13077 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3599
  signal tmp_ivl_1308 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2985
  signal tmp_ivl_13082 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3599
  signal tmp_ivl_13085 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3599
  signal tmp_ivl_13086 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3599
  signal tmp_ivl_1309 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2985
  signal tmp_ivl_13091 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3599
  signal tmp_ivl_13093 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3599
  signal tmp_ivl_13099 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3600
  signal tmp_ivl_131 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2944
  signal tmp_ivl_13101 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3600
  signal tmp_ivl_13102 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3600
  signal tmp_ivl_13107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3600
  signal tmp_ivl_13109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3600
  signal tmp_ivl_13114 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3600
  signal tmp_ivl_13116 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3600
  signal tmp_ivl_13121 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3601
  signal tmp_ivl_13126 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3601
  signal tmp_ivl_13128 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3601
  signal tmp_ivl_13133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3601
  signal tmp_ivl_13135 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3601
  signal tmp_ivl_13137 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3601
  signal tmp_ivl_13139 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3601
  signal tmp_ivl_1314 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2985
  signal tmp_ivl_13144 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3602
  signal tmp_ivl_13149 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3602
  signal tmp_ivl_13151 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3602
  signal tmp_ivl_13156 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3602
  signal tmp_ivl_13158 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3602
  signal tmp_ivl_13164 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3603
  signal tmp_ivl_13166 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3603
  signal tmp_ivl_13167 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3603
  signal tmp_ivl_1317 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2985
  signal tmp_ivl_13172 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3603
  signal tmp_ivl_13175 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3603
  signal tmp_ivl_13176 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3603
  signal tmp_ivl_13181 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3603
  signal tmp_ivl_13183 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3603
  signal tmp_ivl_13189 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3604
  signal tmp_ivl_1319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2985
  signal tmp_ivl_13191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3604
  signal tmp_ivl_13192 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3604
  signal tmp_ivl_13197 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3604
  signal tmp_ivl_13199 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3604
  signal tmp_ivl_1320 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2985
  signal tmp_ivl_13204 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3604
  signal tmp_ivl_13206 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3604
  signal tmp_ivl_13211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3605
  signal tmp_ivl_13216 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3605
  signal tmp_ivl_13218 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3605
  signal tmp_ivl_13223 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3605
  signal tmp_ivl_13225 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3605
  signal tmp_ivl_13227 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3605
  signal tmp_ivl_13229 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3605
  signal tmp_ivl_13234 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3606
  signal tmp_ivl_13239 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3606
  signal tmp_ivl_13241 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3606
  signal tmp_ivl_13246 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3606
  signal tmp_ivl_13248 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3606
  signal tmp_ivl_1325 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2985
  signal tmp_ivl_13253 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3607
  signal tmp_ivl_13258 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3607
  signal tmp_ivl_13260 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3607
  signal tmp_ivl_13265 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3607
  signal tmp_ivl_13267 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3607
  signal tmp_ivl_13269 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3607
  signal tmp_ivl_1327 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2985
  signal tmp_ivl_13271 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3607
  signal tmp_ivl_13277 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3608
  signal tmp_ivl_13278 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3608
  signal tmp_ivl_13283 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3608
  signal tmp_ivl_13286 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3608
  signal tmp_ivl_13288 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3608
  signal tmp_ivl_13289 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3608
  signal tmp_ivl_1329 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2985
  signal tmp_ivl_13294 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3608
  signal tmp_ivl_13296 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3608
  signal tmp_ivl_13302 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3609
  signal tmp_ivl_13303 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3609
  signal tmp_ivl_13308 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3609
  signal tmp_ivl_13311 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3609
  signal tmp_ivl_13313 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3609
  signal tmp_ivl_13314 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3609
  signal tmp_ivl_13319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3609
  signal tmp_ivl_13321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3609
  signal tmp_ivl_13327 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3610
  signal tmp_ivl_13329 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3610
  signal tmp_ivl_13330 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3610
  signal tmp_ivl_13335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3610
  signal tmp_ivl_13337 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3610
  signal tmp_ivl_13342 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3610
  signal tmp_ivl_13344 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3610
  signal tmp_ivl_13349 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3611
  signal tmp_ivl_1335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2986
  signal tmp_ivl_13354 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3611
  signal tmp_ivl_13356 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3611
  signal tmp_ivl_13361 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3611
  signal tmp_ivl_13363 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3611
  signal tmp_ivl_13368 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3612
  signal tmp_ivl_1337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2986
  signal tmp_ivl_13373 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3612
  signal tmp_ivl_13375 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3612
  signal tmp_ivl_1338 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2986
  signal tmp_ivl_13380 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3612
  signal tmp_ivl_13382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3612
  signal tmp_ivl_13388 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3613
  signal tmp_ivl_13389 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3613
  signal tmp_ivl_13394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3613
  signal tmp_ivl_13397 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3613
  signal tmp_ivl_13399 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3613
  signal tmp_ivl_13400 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3613
  signal tmp_ivl_13405 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3613
  signal tmp_ivl_13407 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3613
  signal tmp_ivl_13413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3614
  signal tmp_ivl_13414 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3614
  signal tmp_ivl_13419 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3614
  signal tmp_ivl_13422 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3614
  signal tmp_ivl_13424 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3614
  signal tmp_ivl_13425 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3614
  signal tmp_ivl_1343 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2986
  signal tmp_ivl_13430 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3614
  signal tmp_ivl_13432 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3614
  signal tmp_ivl_13438 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3615
  signal tmp_ivl_13440 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3615
  signal tmp_ivl_13441 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3615
  signal tmp_ivl_13446 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3615
  signal tmp_ivl_13448 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3615
  signal tmp_ivl_13453 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3615
  signal tmp_ivl_13455 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3615
  signal tmp_ivl_1346 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2986
  signal tmp_ivl_13460 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3616
  signal tmp_ivl_13465 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3616
  signal tmp_ivl_13467 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3616
  signal tmp_ivl_13472 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3616
  signal tmp_ivl_13474 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3616
  signal tmp_ivl_13479 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3617
  signal tmp_ivl_1348 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2986
  signal tmp_ivl_13484 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3617
  signal tmp_ivl_13486 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3617
  signal tmp_ivl_1349 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2986
  signal tmp_ivl_13491 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3617
  signal tmp_ivl_13493 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3617
  signal tmp_ivl_13495 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3617
  signal tmp_ivl_13497 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3617
  signal tmp_ivl_13503 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3618
  signal tmp_ivl_13504 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3618
  signal tmp_ivl_13509 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3618
  signal tmp_ivl_13512 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3618
  signal tmp_ivl_13514 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3618
  signal tmp_ivl_13515 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3618
  signal tmp_ivl_13520 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3618
  signal tmp_ivl_13522 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3618
  signal tmp_ivl_13528 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3619
  signal tmp_ivl_13529 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3619
  signal tmp_ivl_13534 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3619
  signal tmp_ivl_13537 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3619
  signal tmp_ivl_13539 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3619
  signal tmp_ivl_1354 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2986
  signal tmp_ivl_13540 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3619
  signal tmp_ivl_13545 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3619
  signal tmp_ivl_13547 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3619
  signal tmp_ivl_13553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3620
  signal tmp_ivl_13555 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3620
  signal tmp_ivl_13556 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3620
  signal tmp_ivl_1356 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2986
  signal tmp_ivl_13561 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3620
  signal tmp_ivl_13563 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3620
  signal tmp_ivl_13568 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3620
  signal tmp_ivl_13570 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3620
  signal tmp_ivl_13575 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3621
  signal tmp_ivl_1358 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2986
  signal tmp_ivl_13580 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3621
  signal tmp_ivl_13582 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3621
  signal tmp_ivl_13587 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3621
  signal tmp_ivl_13589 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3621
  signal tmp_ivl_13595 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3622
  signal tmp_ivl_13596 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3622
  signal tmp_ivl_136 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2944
  signal tmp_ivl_13601 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3622
  signal tmp_ivl_13604 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3622
  signal tmp_ivl_13606 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3622
  signal tmp_ivl_13607 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3622
  signal tmp_ivl_13612 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3622
  signal tmp_ivl_13614 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3622
  signal tmp_ivl_13620 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3623
  signal tmp_ivl_13621 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3623
  signal tmp_ivl_13626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3623
  signal tmp_ivl_13628 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3623
  signal tmp_ivl_13633 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3623
  signal tmp_ivl_13635 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3623
  signal tmp_ivl_1364 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2987
  signal tmp_ivl_13640 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3624
  signal tmp_ivl_13645 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3624
  signal tmp_ivl_13647 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3624
  signal tmp_ivl_13652 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3624
  signal tmp_ivl_13654 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3624
  signal tmp_ivl_13659 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3625
  signal tmp_ivl_1366 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2987
  signal tmp_ivl_13664 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3625
  signal tmp_ivl_13666 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3625
  signal tmp_ivl_1367 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2987
  signal tmp_ivl_13671 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3625
  signal tmp_ivl_13673 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3625
  signal tmp_ivl_13679 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3626
  signal tmp_ivl_13680 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3626
  signal tmp_ivl_13685 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3626
  signal tmp_ivl_13688 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3626
  signal tmp_ivl_13690 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3626
  signal tmp_ivl_13691 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3626
  signal tmp_ivl_13696 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3626
  signal tmp_ivl_13698 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3626
  signal tmp_ivl_13704 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3627
  signal tmp_ivl_13705 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3627
  signal tmp_ivl_13710 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3627
  signal tmp_ivl_13712 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3627
  signal tmp_ivl_13717 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3627
  signal tmp_ivl_13719 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3627
  signal tmp_ivl_1372 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2987
  signal tmp_ivl_13724 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3628
  signal tmp_ivl_13729 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3628
  signal tmp_ivl_13731 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3628
  signal tmp_ivl_13736 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3628
  signal tmp_ivl_13738 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3628
  signal tmp_ivl_13743 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3629
  signal tmp_ivl_13748 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3629
  signal tmp_ivl_1375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2987
  signal tmp_ivl_13750 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3629
  signal tmp_ivl_13755 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3629
  signal tmp_ivl_13757 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3629
  signal tmp_ivl_13759 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3629
  signal tmp_ivl_13761 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3629
  signal tmp_ivl_13766 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3630
  signal tmp_ivl_1377 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2987
  signal tmp_ivl_13771 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3630
  signal tmp_ivl_13773 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3630
  signal tmp_ivl_13778 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3630
  signal tmp_ivl_1378 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2987
  signal tmp_ivl_13780 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3630
  signal tmp_ivl_13786 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3631
  signal tmp_ivl_13788 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3631
  signal tmp_ivl_13789 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3631
  signal tmp_ivl_13794 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3631
  signal tmp_ivl_13797 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3631
  signal tmp_ivl_13798 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3631
  signal tmp_ivl_138 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2944
  signal tmp_ivl_13803 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3631
  signal tmp_ivl_13805 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3631
  signal tmp_ivl_13811 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3632
  signal tmp_ivl_13813 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3632
  signal tmp_ivl_13814 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3632
  signal tmp_ivl_13819 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3632
  signal tmp_ivl_13821 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3632
  signal tmp_ivl_13826 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3632
  signal tmp_ivl_13828 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3632
  signal tmp_ivl_1383 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2987
  signal tmp_ivl_13833 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3633
  signal tmp_ivl_13838 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3633
  signal tmp_ivl_13840 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3633
  signal tmp_ivl_13845 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3633
  signal tmp_ivl_13847 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3633
  signal tmp_ivl_13849 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3633
  signal tmp_ivl_1385 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2987
  signal tmp_ivl_13851 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3633
  signal tmp_ivl_13856 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3634
  signal tmp_ivl_13861 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3634
  signal tmp_ivl_13863 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3634
  signal tmp_ivl_13868 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3634
  signal tmp_ivl_1387 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2987
  signal tmp_ivl_13870 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3634
  signal tmp_ivl_13875 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3635
  signal tmp_ivl_13880 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3635
  signal tmp_ivl_13882 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3635
  signal tmp_ivl_13887 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3635
  signal tmp_ivl_13889 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3635
  signal tmp_ivl_13891 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3635
  signal tmp_ivl_13893 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3635
  signal tmp_ivl_13898 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3636
  signal tmp_ivl_13903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3636
  signal tmp_ivl_13905 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3636
  signal tmp_ivl_13910 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3636
  signal tmp_ivl_13912 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3636
  signal tmp_ivl_13917 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3637
  signal tmp_ivl_13922 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3637
  signal tmp_ivl_13924 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3637
  signal tmp_ivl_13929 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3637
  signal tmp_ivl_1393 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2988
  signal tmp_ivl_13931 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3637
  signal tmp_ivl_13937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3638
  signal tmp_ivl_13938 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3638
  signal tmp_ivl_13943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3638
  signal tmp_ivl_13946 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3638
  signal tmp_ivl_13948 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3638
  signal tmp_ivl_13949 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3638
  signal tmp_ivl_1395 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2988
  signal tmp_ivl_13954 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3638
  signal tmp_ivl_13956 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3638
  signal tmp_ivl_1396 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2988
  signal tmp_ivl_13961 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3639
  signal tmp_ivl_13966 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3639
  signal tmp_ivl_13968 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3639
  signal tmp_ivl_13973 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3639
  signal tmp_ivl_13975 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3639
  signal tmp_ivl_13980 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3640
  signal tmp_ivl_13985 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3640
  signal tmp_ivl_13987 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3640
  signal tmp_ivl_13992 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3640
  signal tmp_ivl_13994 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3640
  signal tmp_ivl_13996 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3640
  signal tmp_ivl_13998 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3640
  signal tmp_ivl_14 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2940
  signal tmp_ivl_140 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2944
  signal tmp_ivl_14004 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3641
  signal tmp_ivl_14005 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3641
  signal tmp_ivl_1401 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2988
  signal tmp_ivl_14010 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3641
  signal tmp_ivl_14013 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3641
  signal tmp_ivl_14015 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3641
  signal tmp_ivl_14016 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3641
  signal tmp_ivl_14021 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3641
  signal tmp_ivl_14023 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3641
  signal tmp_ivl_14029 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3642
  signal tmp_ivl_14031 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3642
  signal tmp_ivl_14032 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3642
  signal tmp_ivl_14037 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3642
  signal tmp_ivl_14039 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3642
  signal tmp_ivl_1404 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2988
  signal tmp_ivl_14044 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3642
  signal tmp_ivl_14046 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3642
  signal tmp_ivl_14051 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3643
  signal tmp_ivl_14056 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3643
  signal tmp_ivl_14058 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3643
  signal tmp_ivl_1406 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2988
  signal tmp_ivl_14063 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3643
  signal tmp_ivl_14065 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3643
  signal tmp_ivl_1407 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2988
  signal tmp_ivl_14070 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3644
  signal tmp_ivl_14075 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3644
  signal tmp_ivl_14077 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3644
  signal tmp_ivl_14082 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3644
  signal tmp_ivl_14084 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3644
  signal tmp_ivl_14090 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3645
  signal tmp_ivl_14091 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3645
  signal tmp_ivl_14096 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3645
  signal tmp_ivl_14099 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3645
  signal tmp_ivl_14101 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3645
  signal tmp_ivl_14102 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3645
  signal tmp_ivl_14107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3645
  signal tmp_ivl_14109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3645
  signal tmp_ivl_14115 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3646
  signal tmp_ivl_14116 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3646
  signal tmp_ivl_1412 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2988
  signal tmp_ivl_14121 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3646
  signal tmp_ivl_14124 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3646
  signal tmp_ivl_14126 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3646
  signal tmp_ivl_14127 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3646
  signal tmp_ivl_14132 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3646
  signal tmp_ivl_14134 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3646
  signal tmp_ivl_1414 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2988
  signal tmp_ivl_14140 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3647
  signal tmp_ivl_14142 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3647
  signal tmp_ivl_14143 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3647
  signal tmp_ivl_14148 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3647
  signal tmp_ivl_14150 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3647
  signal tmp_ivl_14155 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3647
  signal tmp_ivl_14157 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3647
  signal tmp_ivl_1416 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2988
  signal tmp_ivl_14162 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3648
  signal tmp_ivl_14167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3648
  signal tmp_ivl_14169 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3648
  signal tmp_ivl_14174 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3648
  signal tmp_ivl_14176 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3648
  signal tmp_ivl_14181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3649
  signal tmp_ivl_14186 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3649
  signal tmp_ivl_14188 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3649
  signal tmp_ivl_14193 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3649
  signal tmp_ivl_14195 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3649
  signal tmp_ivl_14197 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3649
  signal tmp_ivl_14199 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3649
  signal tmp_ivl_14205 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3650
  signal tmp_ivl_14206 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3650
  signal tmp_ivl_14211 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3650
  signal tmp_ivl_14214 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3650
  signal tmp_ivl_14216 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3650
  signal tmp_ivl_14217 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3650
  signal tmp_ivl_1422 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2989
  signal tmp_ivl_14222 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3650
  signal tmp_ivl_14224 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3650
  signal tmp_ivl_14229 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3651
  signal tmp_ivl_14234 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3651
  signal tmp_ivl_14236 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3651
  signal tmp_ivl_1424 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2989
  signal tmp_ivl_14241 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3651
  signal tmp_ivl_14243 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3651
  signal tmp_ivl_14249 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3652
  signal tmp_ivl_1425 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2989
  signal tmp_ivl_14250 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3652
  signal tmp_ivl_14255 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3652
  signal tmp_ivl_14258 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3652
  signal tmp_ivl_14260 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3652
  signal tmp_ivl_14261 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3652
  signal tmp_ivl_14266 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3652
  signal tmp_ivl_14268 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3652
  signal tmp_ivl_14273 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3653
  signal tmp_ivl_14278 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3653
  signal tmp_ivl_14280 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3653
  signal tmp_ivl_14285 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3653
  signal tmp_ivl_14287 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3653
  signal tmp_ivl_14292 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3654
  signal tmp_ivl_14297 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3654
  signal tmp_ivl_14299 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3654
  signal tmp_ivl_1430 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2989
  signal tmp_ivl_14304 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3654
  signal tmp_ivl_14306 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3654
  signal tmp_ivl_14311 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3655
  signal tmp_ivl_14316 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3655
  signal tmp_ivl_14318 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3655
  signal tmp_ivl_14323 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3655
  signal tmp_ivl_14325 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3655
  signal tmp_ivl_1433 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2989
  signal tmp_ivl_14330 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3656
  signal tmp_ivl_14335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3656
  signal tmp_ivl_14337 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3656
  signal tmp_ivl_14342 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3656
  signal tmp_ivl_14344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3656
  signal tmp_ivl_14346 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3656
  signal tmp_ivl_14348 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3656
  signal tmp_ivl_1435 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2989
  signal tmp_ivl_14354 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3657
  signal tmp_ivl_14355 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3657
  signal tmp_ivl_1436 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2989
  signal tmp_ivl_14360 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3657
  signal tmp_ivl_14363 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3657
  signal tmp_ivl_14365 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3657
  signal tmp_ivl_14366 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3657
  signal tmp_ivl_14371 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3657
  signal tmp_ivl_14373 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3657
  signal tmp_ivl_14379 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3658
  signal tmp_ivl_14381 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3658
  signal tmp_ivl_14382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3658
  signal tmp_ivl_14387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3658
  signal tmp_ivl_14389 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3658
  signal tmp_ivl_14394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3658
  signal tmp_ivl_14396 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3658
  signal tmp_ivl_14401 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3659
  signal tmp_ivl_14406 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3659
  signal tmp_ivl_14408 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3659
  signal tmp_ivl_1441 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2989
  signal tmp_ivl_14413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3659
  signal tmp_ivl_14415 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3659
  signal tmp_ivl_14420 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3660
  signal tmp_ivl_14425 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3660
  signal tmp_ivl_14427 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3660
  signal tmp_ivl_1443 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2989
  signal tmp_ivl_14432 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3660
  signal tmp_ivl_14434 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3660
  signal tmp_ivl_14440 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3661
  signal tmp_ivl_14441 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3661
  signal tmp_ivl_14446 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3661
  signal tmp_ivl_14449 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3661
  signal tmp_ivl_1445 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2989
  signal tmp_ivl_14451 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3661
  signal tmp_ivl_14452 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3661
  signal tmp_ivl_14457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3661
  signal tmp_ivl_14459 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3661
  signal tmp_ivl_14465 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3662
  signal tmp_ivl_14467 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3662
  signal tmp_ivl_14468 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3662
  signal tmp_ivl_14473 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3662
  signal tmp_ivl_14475 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3662
  signal tmp_ivl_14480 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3662
  signal tmp_ivl_14482 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3662
  signal tmp_ivl_14487 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3663
  signal tmp_ivl_14492 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3663
  signal tmp_ivl_14494 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3663
  signal tmp_ivl_14499 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3663
  signal tmp_ivl_14501 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3663
  signal tmp_ivl_14506 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3664
  signal tmp_ivl_1451 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2990
  signal tmp_ivl_14511 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3664
  signal tmp_ivl_14513 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3664
  signal tmp_ivl_14518 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3664
  signal tmp_ivl_14520 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3664
  signal tmp_ivl_14522 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3664
  signal tmp_ivl_14524 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3664
  signal tmp_ivl_14529 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3665
  signal tmp_ivl_1453 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2990
  signal tmp_ivl_14534 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3665
  signal tmp_ivl_14536 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3665
  signal tmp_ivl_1454 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2990
  signal tmp_ivl_14541 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3665
  signal tmp_ivl_14543 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3665
  signal tmp_ivl_14548 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3666
  signal tmp_ivl_14553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3666
  signal tmp_ivl_14555 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3666
  signal tmp_ivl_14560 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3666
  signal tmp_ivl_14562 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3666
  signal tmp_ivl_14564 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3666
  signal tmp_ivl_14566 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3666
  signal tmp_ivl_14572 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3667
  signal tmp_ivl_14573 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3667
  signal tmp_ivl_14578 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3667
  signal tmp_ivl_14581 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3667
  signal tmp_ivl_14583 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3667
  signal tmp_ivl_14584 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3667
  signal tmp_ivl_14589 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3667
  signal tmp_ivl_1459 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2990
  signal tmp_ivl_14591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3667
  signal tmp_ivl_14597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3668
  signal tmp_ivl_14599 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3668
  signal tmp_ivl_146 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2945
  signal tmp_ivl_14600 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3668
  signal tmp_ivl_14605 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3668
  signal tmp_ivl_14608 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3668
  signal tmp_ivl_14609 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3668
  signal tmp_ivl_14614 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3668
  signal tmp_ivl_14616 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3668
  signal tmp_ivl_1462 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2990
  signal tmp_ivl_14621 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3669
  signal tmp_ivl_14626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3669
  signal tmp_ivl_14628 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3669
  signal tmp_ivl_14633 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3669
  signal tmp_ivl_14635 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3669
  signal tmp_ivl_1464 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2990
  signal tmp_ivl_14641 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3670
  signal tmp_ivl_14642 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3670
  signal tmp_ivl_14647 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3670
  signal tmp_ivl_1465 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2990
  signal tmp_ivl_14650 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3670
  signal tmp_ivl_14652 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3670
  signal tmp_ivl_14653 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3670
  signal tmp_ivl_14658 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3670
  signal tmp_ivl_14660 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3670
  signal tmp_ivl_14665 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3671
  signal tmp_ivl_14670 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3671
  signal tmp_ivl_14672 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3671
  signal tmp_ivl_14677 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3671
  signal tmp_ivl_14679 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3671
  signal tmp_ivl_14684 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3672
  signal tmp_ivl_14689 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3672
  signal tmp_ivl_14691 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3672
  signal tmp_ivl_14696 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3672
  signal tmp_ivl_14698 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3672
  signal tmp_ivl_1470 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2990
  signal tmp_ivl_14703 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3673
  signal tmp_ivl_14708 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3673
  signal tmp_ivl_14710 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3673
  signal tmp_ivl_14715 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3673
  signal tmp_ivl_14717 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3673
  signal tmp_ivl_1472 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2990
  signal tmp_ivl_14722 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3674
  signal tmp_ivl_14727 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3674
  signal tmp_ivl_14729 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3674
  signal tmp_ivl_14734 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3674
  signal tmp_ivl_14736 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3674
  signal tmp_ivl_14738 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3674
  signal tmp_ivl_1474 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2990
  signal tmp_ivl_14740 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3674
  signal tmp_ivl_14745 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3675
  signal tmp_ivl_14750 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3675
  signal tmp_ivl_14752 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3675
  signal tmp_ivl_14757 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3675
  signal tmp_ivl_14759 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3675
  signal tmp_ivl_14765 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3676
  signal tmp_ivl_14767 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3676
  signal tmp_ivl_14768 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3676
  signal tmp_ivl_14773 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3676
  signal tmp_ivl_14775 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3676
  signal tmp_ivl_14780 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3676
  signal tmp_ivl_14782 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3676
  signal tmp_ivl_14787 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3677
  signal tmp_ivl_14792 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3677
  signal tmp_ivl_14794 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3677
  signal tmp_ivl_14799 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3677
  signal tmp_ivl_148 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2945
  signal tmp_ivl_1480 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2991
  signal tmp_ivl_14801 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3677
  signal tmp_ivl_14803 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3677
  signal tmp_ivl_14805 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3677
  signal tmp_ivl_14811 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3678
  signal tmp_ivl_14812 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3678
  signal tmp_ivl_14817 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3678
  signal tmp_ivl_1482 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2991
  signal tmp_ivl_14820 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3678
  signal tmp_ivl_14822 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3678
  signal tmp_ivl_14823 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3678
  signal tmp_ivl_14828 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3678
  signal tmp_ivl_1483 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2991
  signal tmp_ivl_14830 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3678
  signal tmp_ivl_14836 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3679
  signal tmp_ivl_14837 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3679
  signal tmp_ivl_14842 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3679
  signal tmp_ivl_14845 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3679
  signal tmp_ivl_14847 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3679
  signal tmp_ivl_14848 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3679
  signal tmp_ivl_14853 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3679
  signal tmp_ivl_14855 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3679
  signal tmp_ivl_14861 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3680
  signal tmp_ivl_14863 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3680
  signal tmp_ivl_14864 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3680
  signal tmp_ivl_14869 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3680
  signal tmp_ivl_14871 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3680
  signal tmp_ivl_14876 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3680
  signal tmp_ivl_14878 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3680
  signal tmp_ivl_1488 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2991
  signal tmp_ivl_14883 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3681
  signal tmp_ivl_14888 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3681
  signal tmp_ivl_14890 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3681
  signal tmp_ivl_14895 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3681
  signal tmp_ivl_14897 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3681
  signal tmp_ivl_149 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2945
  signal tmp_ivl_14903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3682
  signal tmp_ivl_14904 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3682
  signal tmp_ivl_14909 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3682
  signal tmp_ivl_1491 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2991
  signal tmp_ivl_14912 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3682
  signal tmp_ivl_14914 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3682
  signal tmp_ivl_14915 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3682
  signal tmp_ivl_14920 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3682
  signal tmp_ivl_14922 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3682
  signal tmp_ivl_14928 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3683
  signal tmp_ivl_1493 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2991
  signal tmp_ivl_14930 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3683
  signal tmp_ivl_14931 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3683
  signal tmp_ivl_14936 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3683
  signal tmp_ivl_14938 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3683
  signal tmp_ivl_1494 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2991
  signal tmp_ivl_14943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3683
  signal tmp_ivl_14945 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3683
  signal tmp_ivl_14950 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3684
  signal tmp_ivl_14955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3684
  signal tmp_ivl_14957 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3684
  signal tmp_ivl_14962 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3684
  signal tmp_ivl_14964 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3684
  signal tmp_ivl_14969 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3685
  signal tmp_ivl_14974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3685
  signal tmp_ivl_14976 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3685
  signal tmp_ivl_14981 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3685
  signal tmp_ivl_14983 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3685
  signal tmp_ivl_14989 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3686
  signal tmp_ivl_1499 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2991
  signal tmp_ivl_14990 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3686
  signal tmp_ivl_14995 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3686
  signal tmp_ivl_14998 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3686
  signal tmp_ivl_15 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2940
  signal tmp_ivl_15000 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3686
  signal tmp_ivl_15001 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3686
  signal tmp_ivl_15006 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3686
  signal tmp_ivl_15008 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3686
  signal tmp_ivl_1501 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2991
  signal tmp_ivl_15014 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3687
  signal tmp_ivl_15015 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3687
  signal tmp_ivl_15020 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3687
  signal tmp_ivl_15022 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3687
  signal tmp_ivl_15027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3687
  signal tmp_ivl_15029 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3687
  signal tmp_ivl_1503 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2991
  signal tmp_ivl_15034 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3688
  signal tmp_ivl_15039 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3688
  signal tmp_ivl_15041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3688
  signal tmp_ivl_15046 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3688
  signal tmp_ivl_15048 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3688
  signal tmp_ivl_15053 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3689
  signal tmp_ivl_15058 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3689
  signal tmp_ivl_15060 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3689
  signal tmp_ivl_15065 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3689
  signal tmp_ivl_15067 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3689
  signal tmp_ivl_15069 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3689
  signal tmp_ivl_15071 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3689
  signal tmp_ivl_15076 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3690
  signal tmp_ivl_15081 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3690
  signal tmp_ivl_15083 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3690
  signal tmp_ivl_15088 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3690
  signal tmp_ivl_1509 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2992
  signal tmp_ivl_15090 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3690
  signal tmp_ivl_15095 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3691
  signal tmp_ivl_15100 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3691
  signal tmp_ivl_15102 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3691
  signal tmp_ivl_15107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3691
  signal tmp_ivl_15109 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3691
  signal tmp_ivl_1511 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2992
  signal tmp_ivl_15111 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3691
  signal tmp_ivl_15113 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3691
  signal tmp_ivl_15118 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3692
  signal tmp_ivl_1512 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2992
  signal tmp_ivl_15123 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3692
  signal tmp_ivl_15125 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3692
  signal tmp_ivl_15130 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3692
  signal tmp_ivl_15132 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3692
  signal tmp_ivl_15137 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3693
  signal tmp_ivl_15142 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3693
  signal tmp_ivl_15144 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3693
  signal tmp_ivl_15149 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3693
  signal tmp_ivl_15151 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3693
  signal tmp_ivl_15153 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3693
  signal tmp_ivl_15155 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3693
  signal tmp_ivl_15161 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3694
  signal tmp_ivl_15162 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3694
  signal tmp_ivl_15167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3694
  signal tmp_ivl_1517 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2992
  signal tmp_ivl_15170 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3694
  signal tmp_ivl_15172 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3694
  signal tmp_ivl_15173 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3694
  signal tmp_ivl_15178 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3694
  signal tmp_ivl_15180 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3694
  signal tmp_ivl_15185 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3695
  signal tmp_ivl_15190 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3695
  signal tmp_ivl_15192 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3695
  signal tmp_ivl_15197 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3695
  signal tmp_ivl_15199 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3695
  signal tmp_ivl_1520 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2992
  signal tmp_ivl_15204 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3696
  signal tmp_ivl_15209 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3696
  signal tmp_ivl_15211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3696
  signal tmp_ivl_15216 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3696
  signal tmp_ivl_15218 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3696
  signal tmp_ivl_1522 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2992
  signal tmp_ivl_15223 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3697
  signal tmp_ivl_15228 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3697
  signal tmp_ivl_1523 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2992
  signal tmp_ivl_15230 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3697
  signal tmp_ivl_15235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3697
  signal tmp_ivl_15237 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3697
  signal tmp_ivl_15242 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3698
  signal tmp_ivl_15247 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3698
  signal tmp_ivl_15249 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3698
  signal tmp_ivl_15254 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3698
  signal tmp_ivl_15256 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3698
  signal tmp_ivl_15261 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3699
  signal tmp_ivl_15266 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3699
  signal tmp_ivl_15268 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3699
  signal tmp_ivl_15273 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3699
  signal tmp_ivl_15275 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3699
  signal tmp_ivl_15277 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3699
  signal tmp_ivl_15279 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3699
  signal tmp_ivl_1528 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2992
  signal tmp_ivl_15285 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3700
  signal tmp_ivl_15286 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3700
  signal tmp_ivl_15291 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3700
  signal tmp_ivl_15294 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3700
  signal tmp_ivl_15296 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3700
  signal tmp_ivl_15297 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3700
  signal tmp_ivl_1530 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2992
  signal tmp_ivl_15302 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3700
  signal tmp_ivl_15304 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3700
  signal tmp_ivl_15310 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3701
  signal tmp_ivl_15312 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3701
  signal tmp_ivl_15313 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3701
  signal tmp_ivl_15318 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3701
  signal tmp_ivl_1532 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2992
  signal tmp_ivl_15320 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3701
  signal tmp_ivl_15325 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3701
  signal tmp_ivl_15327 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3701
  signal tmp_ivl_15332 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3702
  signal tmp_ivl_15337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3702
  signal tmp_ivl_15339 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3702
  signal tmp_ivl_15344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3702
  signal tmp_ivl_15346 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3702
  signal tmp_ivl_15351 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3703
  signal tmp_ivl_15356 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3703
  signal tmp_ivl_15358 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3703
  signal tmp_ivl_15363 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3703
  signal tmp_ivl_15365 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3703
  signal tmp_ivl_15371 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3704
  signal tmp_ivl_15372 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3704
  signal tmp_ivl_15377 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3704
  signal tmp_ivl_15379 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3704
  signal tmp_ivl_1538 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2993
  signal tmp_ivl_15384 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3704
  signal tmp_ivl_15386 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3704
  signal tmp_ivl_15391 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3705
  signal tmp_ivl_15396 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3705
  signal tmp_ivl_15398 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3705
  signal tmp_ivl_154 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2945
  signal tmp_ivl_1540 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2993
  signal tmp_ivl_15403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3705
  signal tmp_ivl_15405 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3705
  signal tmp_ivl_1541 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2993
  signal tmp_ivl_15410 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3706
  signal tmp_ivl_15415 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3706
  signal tmp_ivl_15417 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3706
  signal tmp_ivl_15422 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3706
  signal tmp_ivl_15424 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3706
  signal tmp_ivl_15426 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3706
  signal tmp_ivl_15428 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3706
  signal tmp_ivl_15433 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3707
  signal tmp_ivl_15438 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3707
  signal tmp_ivl_15440 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3707
  signal tmp_ivl_15445 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3707
  signal tmp_ivl_15447 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3707
  signal tmp_ivl_15452 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3708
  signal tmp_ivl_15457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3708
  signal tmp_ivl_15459 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3708
  signal tmp_ivl_1546 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2993
  signal tmp_ivl_15464 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3708
  signal tmp_ivl_15466 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3708
  signal tmp_ivl_15468 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3708
  signal tmp_ivl_15470 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3708
  signal tmp_ivl_15475 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3709
  signal tmp_ivl_15480 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3709
  signal tmp_ivl_15482 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3709
  signal tmp_ivl_15487 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3709
  signal tmp_ivl_15489 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3709
  signal tmp_ivl_1549 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2993
  signal tmp_ivl_15495 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3710
  signal tmp_ivl_15497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3710
  signal tmp_ivl_15498 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3710
  signal tmp_ivl_15503 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3710
  signal tmp_ivl_15506 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3710
  signal tmp_ivl_15507 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3710
  signal tmp_ivl_1551 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2993
  signal tmp_ivl_15512 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3710
  signal tmp_ivl_15514 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3710
  signal tmp_ivl_1552 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2993
  signal tmp_ivl_15520 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3711
  signal tmp_ivl_15522 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3711
  signal tmp_ivl_15523 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3711
  signal tmp_ivl_15528 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3711
  signal tmp_ivl_15530 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3711
  signal tmp_ivl_15535 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3711
  signal tmp_ivl_15537 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3711
  signal tmp_ivl_15542 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3712
  signal tmp_ivl_15547 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3712
  signal tmp_ivl_15549 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3712
  signal tmp_ivl_15554 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3712
  signal tmp_ivl_15556 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3712
  signal tmp_ivl_15558 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3712
  signal tmp_ivl_15560 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3712
  signal tmp_ivl_15565 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3713
  signal tmp_ivl_1557 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2993
  signal tmp_ivl_15570 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3713
  signal tmp_ivl_15572 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3713
  signal tmp_ivl_15577 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3713
  signal tmp_ivl_15579 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3713
  signal tmp_ivl_15584 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3714
  signal tmp_ivl_15589 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3714
  signal tmp_ivl_1559 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2993
  signal tmp_ivl_15591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3714
  signal tmp_ivl_15596 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3714
  signal tmp_ivl_15598 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3714
  signal tmp_ivl_15600 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3714
  signal tmp_ivl_15602 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3714
  signal tmp_ivl_15607 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3715
  signal tmp_ivl_1561 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2993
  signal tmp_ivl_15612 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3715
  signal tmp_ivl_15614 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3715
  signal tmp_ivl_15619 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3715
  signal tmp_ivl_15621 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3715
  signal tmp_ivl_15626 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3716
  signal tmp_ivl_15631 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3716
  signal tmp_ivl_15633 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3716
  signal tmp_ivl_15638 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3716
  signal tmp_ivl_15640 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3716
  signal tmp_ivl_15642 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3716
  signal tmp_ivl_15644 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3716
  signal tmp_ivl_15649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3717
  signal tmp_ivl_15654 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3717
  signal tmp_ivl_15656 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3717
  signal tmp_ivl_15661 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3717
  signal tmp_ivl_15663 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3717
  signal tmp_ivl_15669 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3718
  signal tmp_ivl_1567 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2994
  signal tmp_ivl_15670 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3718
  signal tmp_ivl_15675 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3718
  signal tmp_ivl_15678 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3718
  signal tmp_ivl_15680 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3718
  signal tmp_ivl_15681 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3718
  signal tmp_ivl_15686 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3718
  signal tmp_ivl_15688 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3718
  signal tmp_ivl_1569 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2994
  signal tmp_ivl_15694 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3719
  signal tmp_ivl_15695 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3719
  signal tmp_ivl_157 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2945
  signal tmp_ivl_1570 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2994
  signal tmp_ivl_15700 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3719
  signal tmp_ivl_15703 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3719
  signal tmp_ivl_15705 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3719
  signal tmp_ivl_15706 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3719
  signal tmp_ivl_15711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3719
  signal tmp_ivl_15713 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3719
  signal tmp_ivl_15719 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3720
  signal tmp_ivl_15721 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3720
  signal tmp_ivl_15722 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3720
  signal tmp_ivl_15727 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3720
  signal tmp_ivl_15729 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3720
  signal tmp_ivl_15734 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3720
  signal tmp_ivl_15736 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3720
  signal tmp_ivl_15741 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3721
  signal tmp_ivl_15746 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3721
  signal tmp_ivl_15748 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3721
  signal tmp_ivl_1575 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2994
  signal tmp_ivl_15753 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3721
  signal tmp_ivl_15755 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3721
  signal tmp_ivl_15760 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3722
  signal tmp_ivl_15765 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3722
  signal tmp_ivl_15767 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3722
  signal tmp_ivl_15772 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3722
  signal tmp_ivl_15774 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3722
  signal tmp_ivl_15776 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3722
  signal tmp_ivl_15778 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3722
  signal tmp_ivl_1578 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2994
  signal tmp_ivl_15783 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3723
  signal tmp_ivl_15788 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3723
  signal tmp_ivl_15790 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3723
  signal tmp_ivl_15795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3723
  signal tmp_ivl_15797 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3723
  signal tmp_ivl_1580 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2994
  signal tmp_ivl_15803 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3724
  signal tmp_ivl_15804 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3724
  signal tmp_ivl_15809 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3724
  signal tmp_ivl_1581 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2994
  signal tmp_ivl_15812 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3724
  signal tmp_ivl_15814 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3724
  signal tmp_ivl_15815 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3724
  signal tmp_ivl_15820 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3724
  signal tmp_ivl_15822 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3724
  signal tmp_ivl_15828 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3725
  signal tmp_ivl_15829 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3725
  signal tmp_ivl_15834 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3725
  signal tmp_ivl_15837 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3725
  signal tmp_ivl_15839 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3725
  signal tmp_ivl_15840 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3725
  signal tmp_ivl_15845 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3725
  signal tmp_ivl_15847 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3725
  signal tmp_ivl_15853 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3726
  signal tmp_ivl_15855 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3726
  signal tmp_ivl_15856 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3726
  signal tmp_ivl_1586 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2994
  signal tmp_ivl_15861 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3726
  signal tmp_ivl_15863 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3726
  signal tmp_ivl_15868 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3726
  signal tmp_ivl_15870 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3726
  signal tmp_ivl_15875 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3727
  signal tmp_ivl_1588 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2994
  signal tmp_ivl_15880 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3727
  signal tmp_ivl_15882 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3727
  signal tmp_ivl_15887 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3727
  signal tmp_ivl_15889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3727
  signal tmp_ivl_15894 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3728
  signal tmp_ivl_15899 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3728
  signal tmp_ivl_159 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2945
  signal tmp_ivl_1590 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2994
  signal tmp_ivl_15901 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3728
  signal tmp_ivl_15906 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3728
  signal tmp_ivl_15908 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3728
  signal tmp_ivl_15910 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3728
  signal tmp_ivl_15912 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3728
  signal tmp_ivl_15917 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3729
  signal tmp_ivl_15922 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3729
  signal tmp_ivl_15924 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3729
  signal tmp_ivl_15929 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3729
  signal tmp_ivl_15931 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3729
  signal tmp_ivl_15937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3730
  signal tmp_ivl_15938 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3730
  signal tmp_ivl_15943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3730
  signal tmp_ivl_15946 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3730
  signal tmp_ivl_15948 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3730
  signal tmp_ivl_15949 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3730
  signal tmp_ivl_15954 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3730
  signal tmp_ivl_15956 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3730
  signal tmp_ivl_1596 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2995
  signal tmp_ivl_15962 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3731
  signal tmp_ivl_15963 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3731
  signal tmp_ivl_15968 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3731
  signal tmp_ivl_15970 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3731
  signal tmp_ivl_15975 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3731
  signal tmp_ivl_15977 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3731
  signal tmp_ivl_1598 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2995
  signal tmp_ivl_15982 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3732
  signal tmp_ivl_15987 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3732
  signal tmp_ivl_15989 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3732
  signal tmp_ivl_1599 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2995
  signal tmp_ivl_15994 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3732
  signal tmp_ivl_15996 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3732
  signal tmp_ivl_160 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2945
  signal tmp_ivl_16001 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3733
  signal tmp_ivl_16006 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3733
  signal tmp_ivl_16008 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3733
  signal tmp_ivl_16013 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3733
  signal tmp_ivl_16015 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3733
  signal tmp_ivl_16017 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3733
  signal tmp_ivl_16019 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3733
  signal tmp_ivl_16024 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3734
  signal tmp_ivl_16029 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3734
  signal tmp_ivl_16031 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3734
  signal tmp_ivl_16036 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3734
  signal tmp_ivl_16038 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3734
  signal tmp_ivl_1604 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2995
  signal tmp_ivl_16043 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3735
  signal tmp_ivl_16048 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3735
  signal tmp_ivl_16050 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3735
  signal tmp_ivl_16055 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3735
  signal tmp_ivl_16057 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3735
  signal tmp_ivl_16059 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3735
  signal tmp_ivl_16061 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3735
  signal tmp_ivl_16066 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3736
  signal tmp_ivl_1607 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2995
  signal tmp_ivl_16071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3736
  signal tmp_ivl_16073 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3736
  signal tmp_ivl_16078 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3736
  signal tmp_ivl_16080 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3736
  signal tmp_ivl_16086 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3737
  signal tmp_ivl_16088 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3737
  signal tmp_ivl_16089 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3737
  signal tmp_ivl_1609 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2995
  signal tmp_ivl_16094 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3737
  signal tmp_ivl_16097 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3737
  signal tmp_ivl_16098 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3737
  signal tmp_ivl_1610 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2995
  signal tmp_ivl_16103 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3737
  signal tmp_ivl_16105 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3737
  signal tmp_ivl_16110 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3738
  signal tmp_ivl_16115 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3738
  signal tmp_ivl_16117 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3738
  signal tmp_ivl_16122 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3738
  signal tmp_ivl_16124 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3738
  signal tmp_ivl_16129 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3739
  signal tmp_ivl_16134 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3739
  signal tmp_ivl_16136 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3739
  signal tmp_ivl_16141 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3739
  signal tmp_ivl_16143 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3739
  signal tmp_ivl_16145 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3739
  signal tmp_ivl_16147 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3739
  signal tmp_ivl_1615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2995
  signal tmp_ivl_16153 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3740
  signal tmp_ivl_16154 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3740
  signal tmp_ivl_16159 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3740
  signal tmp_ivl_16162 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3740
  signal tmp_ivl_16164 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3740
  signal tmp_ivl_16165 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3740
  signal tmp_ivl_1617 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2995
  signal tmp_ivl_16170 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3740
  signal tmp_ivl_16172 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3740
  signal tmp_ivl_16177 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3741
  signal tmp_ivl_16182 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3741
  signal tmp_ivl_16184 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3741
  signal tmp_ivl_16189 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3741
  signal tmp_ivl_1619 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2995
  signal tmp_ivl_16191 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3741
  signal tmp_ivl_16196 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3742
  signal tmp_ivl_16201 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3742
  signal tmp_ivl_16203 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3742
  signal tmp_ivl_16208 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3742
  signal tmp_ivl_16210 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3742
  signal tmp_ivl_16215 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3743
  signal tmp_ivl_16220 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3743
  signal tmp_ivl_16222 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3743
  signal tmp_ivl_16227 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3743
  signal tmp_ivl_16229 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3743
  signal tmp_ivl_16234 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3744
  signal tmp_ivl_16239 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3744
  signal tmp_ivl_16241 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3744
  signal tmp_ivl_16246 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3744
  signal tmp_ivl_16248 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3744
  signal tmp_ivl_1625 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2996
  signal tmp_ivl_16250 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3744
  signal tmp_ivl_16252 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3744
  signal tmp_ivl_16257 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3745
  signal tmp_ivl_16262 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3745
  signal tmp_ivl_16264 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3745
  signal tmp_ivl_16269 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3745
  signal tmp_ivl_1627 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2996
  signal tmp_ivl_16271 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3745
  signal tmp_ivl_16277 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3746
  signal tmp_ivl_16279 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3746
  signal tmp_ivl_1628 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2996
  signal tmp_ivl_16280 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3746
  signal tmp_ivl_16285 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3746
  signal tmp_ivl_16287 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3746
  signal tmp_ivl_16292 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3746
  signal tmp_ivl_16294 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3746
  signal tmp_ivl_16299 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3747
  signal tmp_ivl_16304 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3747
  signal tmp_ivl_16306 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3747
  signal tmp_ivl_16311 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3747
  signal tmp_ivl_16313 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3747
  signal tmp_ivl_16315 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3747
  signal tmp_ivl_16317 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3747
  signal tmp_ivl_16323 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3748
  signal tmp_ivl_16324 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3748
  signal tmp_ivl_16329 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3748
  signal tmp_ivl_1633 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2996
  signal tmp_ivl_16332 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3748
  signal tmp_ivl_16334 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3748
  signal tmp_ivl_16335 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3748
  signal tmp_ivl_16340 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3748
  signal tmp_ivl_16342 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3748
  signal tmp_ivl_16347 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3749
  signal tmp_ivl_16352 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3749
  signal tmp_ivl_16354 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3749
  signal tmp_ivl_16359 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3749
  signal tmp_ivl_1636 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2996
  signal tmp_ivl_16361 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3749
  signal tmp_ivl_16366 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3750
  signal tmp_ivl_16371 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3750
  signal tmp_ivl_16373 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3750
  signal tmp_ivl_16378 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3750
  signal tmp_ivl_1638 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2996
  signal tmp_ivl_16380 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3750
  signal tmp_ivl_16385 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3751
  signal tmp_ivl_1639 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2996
  signal tmp_ivl_16390 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3751
  signal tmp_ivl_16392 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3751
  signal tmp_ivl_16397 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3751
  signal tmp_ivl_16399 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3751
  signal tmp_ivl_16405 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3752
  signal tmp_ivl_16406 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3752
  signal tmp_ivl_16411 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3752
  signal tmp_ivl_16414 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3752
  signal tmp_ivl_16416 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3752
  signal tmp_ivl_16417 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3752
  signal tmp_ivl_16422 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3752
  signal tmp_ivl_16424 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3752
  signal tmp_ivl_16429 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3753
  signal tmp_ivl_16434 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3753
  signal tmp_ivl_16436 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3753
  signal tmp_ivl_1644 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2996
  signal tmp_ivl_16441 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3753
  signal tmp_ivl_16443 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3753
  signal tmp_ivl_16448 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3754
  signal tmp_ivl_16453 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3754
  signal tmp_ivl_16455 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3754
  signal tmp_ivl_1646 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2996
  signal tmp_ivl_16460 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3754
  signal tmp_ivl_16462 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3754
  signal tmp_ivl_16464 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3754
  signal tmp_ivl_16466 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3754
  signal tmp_ivl_16471 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3755
  signal tmp_ivl_16476 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3755
  signal tmp_ivl_16478 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3755
  signal tmp_ivl_1648 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2996
  signal tmp_ivl_16483 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3755
  signal tmp_ivl_16485 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3755
  signal tmp_ivl_16491 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3756
  signal tmp_ivl_16492 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3756
  signal tmp_ivl_16497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3756
  signal tmp_ivl_165 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2945
  signal tmp_ivl_16500 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3756
  signal tmp_ivl_16502 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3756
  signal tmp_ivl_16503 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3756
  signal tmp_ivl_16508 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3756
  signal tmp_ivl_16510 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3756
  signal tmp_ivl_16516 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3757
  signal tmp_ivl_16518 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3757
  signal tmp_ivl_16519 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3757
  signal tmp_ivl_16524 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3757
  signal tmp_ivl_16526 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3757
  signal tmp_ivl_16531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3757
  signal tmp_ivl_16533 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3757
  signal tmp_ivl_16538 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3758
  signal tmp_ivl_1654 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2997
  signal tmp_ivl_16543 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3758
  signal tmp_ivl_16545 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3758
  signal tmp_ivl_16550 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3758
  signal tmp_ivl_16552 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3758
  signal tmp_ivl_16557 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3759
  signal tmp_ivl_1656 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2997
  signal tmp_ivl_16562 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3759
  signal tmp_ivl_16564 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3759
  signal tmp_ivl_16569 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3759
  signal tmp_ivl_1657 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2997
  signal tmp_ivl_16571 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3759
  signal tmp_ivl_16573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3759
  signal tmp_ivl_16575 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3759
  signal tmp_ivl_16581 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3760
  signal tmp_ivl_16582 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3760
  signal tmp_ivl_16587 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3760
  signal tmp_ivl_16590 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3760
  signal tmp_ivl_16592 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3760
  signal tmp_ivl_16593 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3760
  signal tmp_ivl_16598 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3760
  signal tmp_ivl_16600 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3760
  signal tmp_ivl_16605 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3761
  signal tmp_ivl_16610 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3761
  signal tmp_ivl_16612 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3761
  signal tmp_ivl_16617 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3761
  signal tmp_ivl_16619 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3761
  signal tmp_ivl_1662 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2997
  signal tmp_ivl_16624 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3762
  signal tmp_ivl_16629 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3762
  signal tmp_ivl_16631 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3762
  signal tmp_ivl_16636 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3762
  signal tmp_ivl_16638 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3762
  signal tmp_ivl_16643 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3763
  signal tmp_ivl_16648 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3763
  signal tmp_ivl_1665 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2997
  signal tmp_ivl_16650 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3763
  signal tmp_ivl_16655 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3763
  signal tmp_ivl_16657 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3763
  signal tmp_ivl_16662 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3764
  signal tmp_ivl_16667 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3764
  signal tmp_ivl_16669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3764
  signal tmp_ivl_1667 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2997
  signal tmp_ivl_16674 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3764
  signal tmp_ivl_16676 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3764
  signal tmp_ivl_1668 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2997
  signal tmp_ivl_16681 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3765
  signal tmp_ivl_16686 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3765
  signal tmp_ivl_16688 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3765
  signal tmp_ivl_16693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3765
  signal tmp_ivl_16695 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3765
  signal tmp_ivl_16697 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3765
  signal tmp_ivl_16699 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3765
  signal tmp_ivl_167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2945
  signal tmp_ivl_16705 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3766
  signal tmp_ivl_16706 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3766
  signal tmp_ivl_16711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3766
  signal tmp_ivl_16714 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3766
  signal tmp_ivl_16716 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3766
  signal tmp_ivl_16717 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3766
  signal tmp_ivl_16722 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3766
  signal tmp_ivl_16724 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3766
  signal tmp_ivl_1673 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2997
  signal tmp_ivl_16730 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3767
  signal tmp_ivl_16732 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3767
  signal tmp_ivl_16733 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3767
  signal tmp_ivl_16738 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3767
  signal tmp_ivl_16740 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3767
  signal tmp_ivl_16745 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3767
  signal tmp_ivl_16747 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3767
  signal tmp_ivl_1675 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2997
  signal tmp_ivl_16752 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3768
  signal tmp_ivl_16757 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3768
  signal tmp_ivl_16759 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3768
  signal tmp_ivl_16764 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3768
  signal tmp_ivl_16766 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3768
  signal tmp_ivl_1677 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2997
  signal tmp_ivl_16771 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3769
  signal tmp_ivl_16776 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3769
  signal tmp_ivl_16778 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3769
  signal tmp_ivl_16783 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3769
  signal tmp_ivl_16785 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3769
  signal tmp_ivl_16791 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3770
  signal tmp_ivl_16792 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3770
  signal tmp_ivl_16797 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3770
  signal tmp_ivl_16800 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3770
  signal tmp_ivl_16802 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3770
  signal tmp_ivl_16803 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3770
  signal tmp_ivl_16808 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3770
  signal tmp_ivl_16810 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3770
  signal tmp_ivl_16816 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3771
  signal tmp_ivl_16818 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3771
  signal tmp_ivl_16819 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3771
  signal tmp_ivl_16824 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3771
  signal tmp_ivl_16826 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3771
  signal tmp_ivl_1683 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2998
  signal tmp_ivl_16831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3771
  signal tmp_ivl_16833 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3771
  signal tmp_ivl_16838 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3772
  signal tmp_ivl_16843 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3772
  signal tmp_ivl_16845 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3772
  signal tmp_ivl_1685 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2998
  signal tmp_ivl_16850 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3772
  signal tmp_ivl_16852 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3772
  signal tmp_ivl_16857 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3773
  signal tmp_ivl_1686 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2998
  signal tmp_ivl_16862 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3773
  signal tmp_ivl_16864 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3773
  signal tmp_ivl_16869 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3773
  signal tmp_ivl_16871 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3773
  signal tmp_ivl_16873 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3773
  signal tmp_ivl_16875 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3773
  signal tmp_ivl_16880 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3774
  signal tmp_ivl_16885 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3774
  signal tmp_ivl_16887 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3774
  signal tmp_ivl_16892 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3774
  signal tmp_ivl_16894 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3774
  signal tmp_ivl_16899 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3775
  signal tmp_ivl_169 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2945
  signal tmp_ivl_16904 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3775
  signal tmp_ivl_16906 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3775
  signal tmp_ivl_1691 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2998
  signal tmp_ivl_16911 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3775
  signal tmp_ivl_16913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3775
  signal tmp_ivl_16915 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3775
  signal tmp_ivl_16917 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3775
  signal tmp_ivl_16922 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3776
  signal tmp_ivl_16927 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3776
  signal tmp_ivl_16929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3776
  signal tmp_ivl_16934 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3776
  signal tmp_ivl_16936 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3776
  signal tmp_ivl_1694 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2998
  signal tmp_ivl_16942 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3777
  signal tmp_ivl_16944 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3777
  signal tmp_ivl_16945 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3777
  signal tmp_ivl_16950 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3777
  signal tmp_ivl_16953 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3777
  signal tmp_ivl_16954 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3777
  signal tmp_ivl_16959 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3777
  signal tmp_ivl_1696 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2998
  signal tmp_ivl_16961 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3777
  signal tmp_ivl_16967 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3778
  signal tmp_ivl_16969 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3778
  signal tmp_ivl_1697 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2998
  signal tmp_ivl_16970 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3778
  signal tmp_ivl_16975 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3778
  signal tmp_ivl_16977 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3778
  signal tmp_ivl_16982 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3778
  signal tmp_ivl_16984 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3778
  signal tmp_ivl_16989 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3779
  signal tmp_ivl_16994 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3779
  signal tmp_ivl_16996 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3779
  signal tmp_ivl_17001 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3779
  signal tmp_ivl_17003 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3779
  signal tmp_ivl_17005 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3779
  signal tmp_ivl_17007 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3779
  signal tmp_ivl_17012 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3780
  signal tmp_ivl_17017 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3780
  signal tmp_ivl_17019 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3780
  signal tmp_ivl_1702 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2998
  signal tmp_ivl_17024 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3780
  signal tmp_ivl_17026 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3780
  signal tmp_ivl_17031 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3781
  signal tmp_ivl_17036 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3781
  signal tmp_ivl_17038 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3781
  signal tmp_ivl_1704 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2998
  signal tmp_ivl_17043 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3781
  signal tmp_ivl_17045 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3781
  signal tmp_ivl_17047 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3781
  signal tmp_ivl_17049 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3781
  signal tmp_ivl_17054 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3782
  signal tmp_ivl_17059 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3782
  signal tmp_ivl_1706 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2998
  signal tmp_ivl_17061 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3782
  signal tmp_ivl_17066 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3782
  signal tmp_ivl_17068 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3782
  signal tmp_ivl_17073 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3783
  signal tmp_ivl_17078 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3783
  signal tmp_ivl_17080 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3783
  signal tmp_ivl_17085 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3783
  signal tmp_ivl_17087 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3783
  signal tmp_ivl_17089 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3783
  signal tmp_ivl_17091 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3783
  signal tmp_ivl_17096 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3784
  signal tmp_ivl_17101 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3784
  signal tmp_ivl_17103 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3784
  signal tmp_ivl_17108 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3784
  signal tmp_ivl_17110 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3784
  signal tmp_ivl_17116 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3785
  signal tmp_ivl_17117 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3785
  signal tmp_ivl_1712 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2999
  signal tmp_ivl_17122 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3785
  signal tmp_ivl_17125 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3785
  signal tmp_ivl_17127 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3785
  signal tmp_ivl_17128 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3785
  signal tmp_ivl_17133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3785
  signal tmp_ivl_17135 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3785
  signal tmp_ivl_1714 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2999
  signal tmp_ivl_17141 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3786
  signal tmp_ivl_17142 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3786
  signal tmp_ivl_17147 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3786
  signal tmp_ivl_1715 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2999
  signal tmp_ivl_17150 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3786
  signal tmp_ivl_17152 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3786
  signal tmp_ivl_17153 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3786
  signal tmp_ivl_17158 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3786
  signal tmp_ivl_17160 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3786
  signal tmp_ivl_17166 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3787
  signal tmp_ivl_17168 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3787
  signal tmp_ivl_17169 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3787
  signal tmp_ivl_17174 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3787
  signal tmp_ivl_17176 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3787
  signal tmp_ivl_17181 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3787
  signal tmp_ivl_17183 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3787
  signal tmp_ivl_17188 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3788
  signal tmp_ivl_17193 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3788
  signal tmp_ivl_17195 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3788
  signal tmp_ivl_1720 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2999
  signal tmp_ivl_17200 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3788
  signal tmp_ivl_17202 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3788
  signal tmp_ivl_17207 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3789
  signal tmp_ivl_17212 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3789
  signal tmp_ivl_17214 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3789
  signal tmp_ivl_17219 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3789
  signal tmp_ivl_17221 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3789
  signal tmp_ivl_17223 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3789
  signal tmp_ivl_17225 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3789
  signal tmp_ivl_1723 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2999
  signal tmp_ivl_17230 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3790
  signal tmp_ivl_17235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3790
  signal tmp_ivl_17237 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3790
  signal tmp_ivl_17242 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3790
  signal tmp_ivl_17244 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3790
  signal tmp_ivl_1725 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2999
  signal tmp_ivl_17250 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3791
  signal tmp_ivl_17251 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3791
  signal tmp_ivl_17256 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3791
  signal tmp_ivl_17259 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3791
  signal tmp_ivl_1726 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2999
  signal tmp_ivl_17261 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3791
  signal tmp_ivl_17262 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3791
  signal tmp_ivl_17267 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3791
  signal tmp_ivl_17269 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3791
  signal tmp_ivl_17275 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3792
  signal tmp_ivl_17276 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3792
  signal tmp_ivl_17281 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3792
  signal tmp_ivl_17283 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3792
  signal tmp_ivl_17288 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3792
  signal tmp_ivl_17290 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3792
  signal tmp_ivl_17295 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3793
  signal tmp_ivl_17300 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3793
  signal tmp_ivl_17302 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3793
  signal tmp_ivl_17307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3793
  signal tmp_ivl_17309 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3793
  signal tmp_ivl_1731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2999
  signal tmp_ivl_17314 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3794
  signal tmp_ivl_17319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3794
  signal tmp_ivl_17321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3794
  signal tmp_ivl_17326 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3794
  signal tmp_ivl_17328 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3794
  signal tmp_ivl_1733 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2999
  signal tmp_ivl_17330 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3794
  signal tmp_ivl_17332 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3794
  signal tmp_ivl_17337 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3795
  signal tmp_ivl_17342 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3795
  signal tmp_ivl_17344 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3795
  signal tmp_ivl_17349 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3795
  signal tmp_ivl_1735 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2999
  signal tmp_ivl_17351 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3795
  signal tmp_ivl_17356 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3796
  signal tmp_ivl_17361 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3796
  signal tmp_ivl_17363 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3796
  signal tmp_ivl_17368 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3796
  signal tmp_ivl_17370 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3796
  signal tmp_ivl_17372 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3796
  signal tmp_ivl_17374 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3796
  signal tmp_ivl_17380 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3797
  signal tmp_ivl_17381 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3797
  signal tmp_ivl_17386 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3797
  signal tmp_ivl_17389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3797
  signal tmp_ivl_17391 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3797
  signal tmp_ivl_17392 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3797
  signal tmp_ivl_17397 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3797
  signal tmp_ivl_17399 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3797
  signal tmp_ivl_17404 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3798
  signal tmp_ivl_17409 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3798
  signal tmp_ivl_1741 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3000
  signal tmp_ivl_17411 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3798
  signal tmp_ivl_17416 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3798
  signal tmp_ivl_17418 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3798
  signal tmp_ivl_17423 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3799
  signal tmp_ivl_17428 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3799
  signal tmp_ivl_1743 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3000
  signal tmp_ivl_17430 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3799
  signal tmp_ivl_17435 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3799
  signal tmp_ivl_17437 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3799
  signal tmp_ivl_1744 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3000
  signal tmp_ivl_17442 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3800
  signal tmp_ivl_17447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3800
  signal tmp_ivl_17449 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3800
  signal tmp_ivl_17454 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3800
  signal tmp_ivl_17456 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3800
  signal tmp_ivl_17461 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3801
  signal tmp_ivl_17466 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3801
  signal tmp_ivl_17468 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3801
  signal tmp_ivl_17473 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3801
  signal tmp_ivl_17475 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3801
  signal tmp_ivl_17477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3801
  signal tmp_ivl_17479 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3801
  signal tmp_ivl_17484 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3802
  signal tmp_ivl_17489 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3802
  signal tmp_ivl_1749 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3000
  signal tmp_ivl_17491 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3802
  signal tmp_ivl_17496 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3802
  signal tmp_ivl_17498 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3802
  signal tmp_ivl_175 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2946
  signal tmp_ivl_17504 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3803
  signal tmp_ivl_17505 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3803
  signal tmp_ivl_17510 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3803
  signal tmp_ivl_17513 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3803
  signal tmp_ivl_17515 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3803
  signal tmp_ivl_17516 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3803
  signal tmp_ivl_1752 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3000
  signal tmp_ivl_17521 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3803
  signal tmp_ivl_17523 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3803
  signal tmp_ivl_17529 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3804
  signal tmp_ivl_17531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3804
  signal tmp_ivl_17532 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3804
  signal tmp_ivl_17537 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3804
  signal tmp_ivl_17539 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3804
  signal tmp_ivl_1754 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3000
  signal tmp_ivl_17544 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3804
  signal tmp_ivl_17546 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3804
  signal tmp_ivl_1755 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3000
  signal tmp_ivl_17551 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3805
  signal tmp_ivl_17556 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3805
  signal tmp_ivl_17558 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3805
  signal tmp_ivl_17563 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3805
  signal tmp_ivl_17565 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3805
  signal tmp_ivl_17570 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3806
  signal tmp_ivl_17575 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3806
  signal tmp_ivl_17577 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3806
  signal tmp_ivl_17582 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3806
  signal tmp_ivl_17584 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3806
  signal tmp_ivl_17586 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3806
  signal tmp_ivl_17588 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3806
  signal tmp_ivl_17593 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3807
  signal tmp_ivl_17598 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3807
  signal tmp_ivl_1760 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3000
  signal tmp_ivl_17600 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3807
  signal tmp_ivl_17605 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3807
  signal tmp_ivl_17607 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3807
  signal tmp_ivl_17613 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3808
  signal tmp_ivl_17615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3808
  signal tmp_ivl_17616 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3808
  signal tmp_ivl_1762 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3000
  signal tmp_ivl_17621 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3808
  signal tmp_ivl_17624 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3808
  signal tmp_ivl_17625 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3808
  signal tmp_ivl_17630 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3808
  signal tmp_ivl_17632 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3808
  signal tmp_ivl_17637 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3809
  signal tmp_ivl_1764 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3000
  signal tmp_ivl_17642 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3809
  signal tmp_ivl_17644 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3809
  signal tmp_ivl_17649 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3809
  signal tmp_ivl_17651 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3809
  signal tmp_ivl_17656 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3810
  signal tmp_ivl_17661 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3810
  signal tmp_ivl_17663 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3810
  signal tmp_ivl_17668 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3810
  signal tmp_ivl_17670 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3810
  signal tmp_ivl_17672 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3810
  signal tmp_ivl_17674 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3810
  signal tmp_ivl_17679 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3811
  signal tmp_ivl_17684 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3811
  signal tmp_ivl_17686 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3811
  signal tmp_ivl_17691 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3811
  signal tmp_ivl_17693 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3811
  signal tmp_ivl_17698 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3812
  signal tmp_ivl_177 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2946
  signal tmp_ivl_1770 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3001
  signal tmp_ivl_17703 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3812
  signal tmp_ivl_17705 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3812
  signal tmp_ivl_17710 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3812
  signal tmp_ivl_17712 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3812
  signal tmp_ivl_17714 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3812
  signal tmp_ivl_17716 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3812
  signal tmp_ivl_1772 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3001
  signal tmp_ivl_17721 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3813
  signal tmp_ivl_17726 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3813
  signal tmp_ivl_17728 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3813
  signal tmp_ivl_1773 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3001
  signal tmp_ivl_17733 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3813
  signal tmp_ivl_17735 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3813
  signal tmp_ivl_17741 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3814
  signal tmp_ivl_17743 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3814
  signal tmp_ivl_17744 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3814
  signal tmp_ivl_17749 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3814
  signal tmp_ivl_17751 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3814
  signal tmp_ivl_17756 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3814
  signal tmp_ivl_17758 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3814
  signal tmp_ivl_17763 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3815
  signal tmp_ivl_17768 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3815
  signal tmp_ivl_17770 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3815
  signal tmp_ivl_17775 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3815
  signal tmp_ivl_17777 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3815
  signal tmp_ivl_17779 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3815
  signal tmp_ivl_1778 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3001
  signal tmp_ivl_17781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3815
  signal tmp_ivl_17786 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3816
  signal tmp_ivl_17791 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3816
  signal tmp_ivl_17793 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3816
  signal tmp_ivl_17798 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3816
  signal tmp_ivl_178 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2946
  signal tmp_ivl_17800 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3816
  signal tmp_ivl_17806 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3817
  signal tmp_ivl_17807 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3817
  signal tmp_ivl_1781 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3001
  signal tmp_ivl_17812 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3817
  signal tmp_ivl_17815 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3817
  signal tmp_ivl_17817 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3817
  signal tmp_ivl_17818 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3817
  signal tmp_ivl_17823 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3817
  signal tmp_ivl_17825 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3817
  signal tmp_ivl_1783 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3001
  signal tmp_ivl_17831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3818
  signal tmp_ivl_17832 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3818
  signal tmp_ivl_17837 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3818
  signal tmp_ivl_1784 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3001
  signal tmp_ivl_17840 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3818
  signal tmp_ivl_17842 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3818
  signal tmp_ivl_17843 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3818
  signal tmp_ivl_17848 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3818
  signal tmp_ivl_17850 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3818
  signal tmp_ivl_17856 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3819
  signal tmp_ivl_17858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3819
  signal tmp_ivl_17859 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3819
  signal tmp_ivl_17864 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3819
  signal tmp_ivl_17866 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3819
  signal tmp_ivl_17871 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3819
  signal tmp_ivl_17873 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3819
  signal tmp_ivl_17878 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3820
  signal tmp_ivl_17883 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3820
  signal tmp_ivl_17885 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3820
  signal tmp_ivl_1789 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3001
  signal tmp_ivl_17890 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3820
  signal tmp_ivl_17892 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3820
  signal tmp_ivl_17897 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3821
  signal tmp_ivl_17902 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3821
  signal tmp_ivl_17904 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3821
  signal tmp_ivl_17909 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3821
  signal tmp_ivl_1791 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3001
  signal tmp_ivl_17911 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3821
  signal tmp_ivl_17913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3821
  signal tmp_ivl_17915 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3821
  signal tmp_ivl_17920 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3822
  signal tmp_ivl_17925 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3822
  signal tmp_ivl_17927 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3822
  signal tmp_ivl_1793 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3001
  signal tmp_ivl_17932 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3822
  signal tmp_ivl_17934 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3822
  signal tmp_ivl_17940 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3823
  signal tmp_ivl_17941 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3823
  signal tmp_ivl_17946 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3823
  signal tmp_ivl_17948 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3823
  signal tmp_ivl_17953 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3823
  signal tmp_ivl_17955 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3823
  signal tmp_ivl_17960 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3824
  signal tmp_ivl_17965 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3824
  signal tmp_ivl_17967 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3824
  signal tmp_ivl_17972 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3824
  signal tmp_ivl_17974 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3824
  signal tmp_ivl_17979 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3825
  signal tmp_ivl_17984 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3825
  signal tmp_ivl_17986 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3825
  signal tmp_ivl_1799 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3002
  signal tmp_ivl_17991 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3825
  signal tmp_ivl_17993 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3825
  signal tmp_ivl_17995 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3825
  signal tmp_ivl_17997 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3825
  signal tmp_ivl_18003 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3826
  signal tmp_ivl_18004 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3826
  signal tmp_ivl_18009 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3826
  signal tmp_ivl_1801 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3002
  signal tmp_ivl_18012 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3826
  signal tmp_ivl_18014 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3826
  signal tmp_ivl_18015 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3826
  signal tmp_ivl_1802 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3002
  signal tmp_ivl_18020 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3826
  signal tmp_ivl_18022 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3826
  signal tmp_ivl_18027 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3827
  signal tmp_ivl_18032 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3827
  signal tmp_ivl_18034 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3827
  signal tmp_ivl_18039 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3827
  signal tmp_ivl_18041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3827
  signal tmp_ivl_18046 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3828
  signal tmp_ivl_18051 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3828
  signal tmp_ivl_18053 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3828
  signal tmp_ivl_18058 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3828
  signal tmp_ivl_18060 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3828
  signal tmp_ivl_18065 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3829
  signal tmp_ivl_1807 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3002
  signal tmp_ivl_18070 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3829
  signal tmp_ivl_18072 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3829
  signal tmp_ivl_18077 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3829
  signal tmp_ivl_18079 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3829
  signal tmp_ivl_18084 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3830
  signal tmp_ivl_18089 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3830
  signal tmp_ivl_18091 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3830
  signal tmp_ivl_18096 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3830
  signal tmp_ivl_18098 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3830
  signal tmp_ivl_1810 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3002
  signal tmp_ivl_18100 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3830
  signal tmp_ivl_18102 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3830
  signal tmp_ivl_18107 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3831
  signal tmp_ivl_18112 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3831
  signal tmp_ivl_18114 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3831
  signal tmp_ivl_18119 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3831
  signal tmp_ivl_1812 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3002
  signal tmp_ivl_18121 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3831
  signal tmp_ivl_18127 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3832
  signal tmp_ivl_18128 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3832
  signal tmp_ivl_1813 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3002
  signal tmp_ivl_18133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3832
  signal tmp_ivl_18136 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3832
  signal tmp_ivl_18138 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3832
  signal tmp_ivl_18139 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3832
  signal tmp_ivl_18144 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3832
  signal tmp_ivl_18146 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3832
  signal tmp_ivl_18152 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3833
  signal tmp_ivl_18154 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3833
  signal tmp_ivl_18155 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3833
  signal tmp_ivl_18160 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3833
  signal tmp_ivl_18162 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3833
  signal tmp_ivl_18167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3833
  signal tmp_ivl_18169 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3833
  signal tmp_ivl_18174 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3834
  signal tmp_ivl_18179 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3834
  signal tmp_ivl_1818 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3002
  signal tmp_ivl_18181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3834
  signal tmp_ivl_18186 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3834
  signal tmp_ivl_18188 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3834
  signal tmp_ivl_18193 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3835
  signal tmp_ivl_18198 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3835
  signal tmp_ivl_1820 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3002
  signal tmp_ivl_18200 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3835
  signal tmp_ivl_18205 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3835
  signal tmp_ivl_18207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3835
  signal tmp_ivl_18209 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3835
  signal tmp_ivl_18211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3835
  signal tmp_ivl_18216 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3836
  signal tmp_ivl_1822 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3002
  signal tmp_ivl_18221 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3836
  signal tmp_ivl_18223 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3836
  signal tmp_ivl_18228 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3836
  signal tmp_ivl_18230 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3836
  signal tmp_ivl_18236 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3837
  signal tmp_ivl_18238 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3837
  signal tmp_ivl_18239 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3837
  signal tmp_ivl_18244 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3837
  signal tmp_ivl_18247 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3837
  signal tmp_ivl_18248 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3837
  signal tmp_ivl_18253 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3837
  signal tmp_ivl_18255 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3837
  signal tmp_ivl_18261 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3838
  signal tmp_ivl_18263 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3838
  signal tmp_ivl_18264 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3838
  signal tmp_ivl_18269 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3838
  signal tmp_ivl_18271 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3838
  signal tmp_ivl_18276 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3838
  signal tmp_ivl_18278 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3838
  signal tmp_ivl_1828 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3003
  signal tmp_ivl_18283 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3839
  signal tmp_ivl_18288 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3839
  signal tmp_ivl_18290 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3839
  signal tmp_ivl_18295 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3839
  signal tmp_ivl_18297 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3839
  signal tmp_ivl_18299 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3839
  signal tmp_ivl_183 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2946
  signal tmp_ivl_1830 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3003
  signal tmp_ivl_18301 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3839
  signal tmp_ivl_18306 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3840
  signal tmp_ivl_1831 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3003
  signal tmp_ivl_18311 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3840
  signal tmp_ivl_18313 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3840
  signal tmp_ivl_18318 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3840
  signal tmp_ivl_18320 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3840
  signal tmp_ivl_18325 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3841
  signal tmp_ivl_18330 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3841
  signal tmp_ivl_18332 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3841
  signal tmp_ivl_18337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3841
  signal tmp_ivl_18339 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3841
  signal tmp_ivl_18341 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3841
  signal tmp_ivl_18343 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3841
  signal tmp_ivl_18348 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3842
  signal tmp_ivl_18353 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3842
  signal tmp_ivl_18355 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3842
  signal tmp_ivl_1836 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3003
  signal tmp_ivl_18360 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3842
  signal tmp_ivl_18362 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3842
  signal tmp_ivl_18367 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3843
  signal tmp_ivl_18372 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3843
  signal tmp_ivl_18374 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3843
  signal tmp_ivl_18379 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3843
  signal tmp_ivl_18381 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3843
  signal tmp_ivl_18383 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3843
  signal tmp_ivl_18385 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3843
  signal tmp_ivl_1839 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3003
  signal tmp_ivl_18391 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3844
  signal tmp_ivl_18392 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3844
  signal tmp_ivl_18397 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3844
  signal tmp_ivl_18400 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3844
  signal tmp_ivl_18402 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3844
  signal tmp_ivl_18403 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3844
  signal tmp_ivl_18408 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3844
  signal tmp_ivl_1841 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3003
  signal tmp_ivl_18410 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3844
  signal tmp_ivl_18415 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3845
  signal tmp_ivl_1842 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3003
  signal tmp_ivl_18420 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3845
  signal tmp_ivl_18422 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3845
  signal tmp_ivl_18427 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3845
  signal tmp_ivl_18429 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3845
  signal tmp_ivl_18434 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3846
  signal tmp_ivl_18439 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3846
  signal tmp_ivl_18441 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3846
  signal tmp_ivl_18446 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3846
  signal tmp_ivl_18448 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3846
  signal tmp_ivl_18453 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3847
  signal tmp_ivl_18458 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3847
  signal tmp_ivl_18460 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3847
  signal tmp_ivl_18465 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3847
  signal tmp_ivl_18467 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3847
  signal tmp_ivl_1847 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3003
  signal tmp_ivl_18472 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3848
  signal tmp_ivl_18477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3848
  signal tmp_ivl_18479 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3848
  signal tmp_ivl_18484 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3848
  signal tmp_ivl_18486 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3848
  signal tmp_ivl_1849 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3003
  signal tmp_ivl_18491 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3849
  signal tmp_ivl_18496 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3849
  signal tmp_ivl_18498 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3849
  signal tmp_ivl_18503 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3849
  signal tmp_ivl_18505 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3849
  signal tmp_ivl_18507 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3849
  signal tmp_ivl_18509 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3849
  signal tmp_ivl_1851 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3003
  signal tmp_ivl_18514 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3850
  signal tmp_ivl_18519 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3850
  signal tmp_ivl_18521 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3850
  signal tmp_ivl_18526 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3850
  signal tmp_ivl_18528 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3850
  signal tmp_ivl_18534 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3851
  signal tmp_ivl_18535 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3851
  signal tmp_ivl_18540 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3851
  signal tmp_ivl_18543 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3851
  signal tmp_ivl_18545 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3851
  signal tmp_ivl_18546 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3851
  signal tmp_ivl_18551 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3851
  signal tmp_ivl_18553 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3851
  signal tmp_ivl_18559 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3852
  signal tmp_ivl_18561 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3852
  signal tmp_ivl_18562 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3852
  signal tmp_ivl_18567 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3852
  signal tmp_ivl_18569 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3852
  signal tmp_ivl_1857 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3004
  signal tmp_ivl_18574 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3852
  signal tmp_ivl_18576 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3852
  signal tmp_ivl_18581 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3853
  signal tmp_ivl_18586 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3853
  signal tmp_ivl_18588 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3853
  signal tmp_ivl_1859 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3004
  signal tmp_ivl_18593 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3853
  signal tmp_ivl_18595 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3853
  signal tmp_ivl_186 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2946
  signal tmp_ivl_1860 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3004
  signal tmp_ivl_18600 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3854
  signal tmp_ivl_18605 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3854
  signal tmp_ivl_18607 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3854
  signal tmp_ivl_18612 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3854
  signal tmp_ivl_18614 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3854
  signal tmp_ivl_18616 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3854
  signal tmp_ivl_18618 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3854
  signal tmp_ivl_18623 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3855
  signal tmp_ivl_18628 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3855
  signal tmp_ivl_18630 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3855
  signal tmp_ivl_18635 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3855
  signal tmp_ivl_18637 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3855
  signal tmp_ivl_18643 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3856
  signal tmp_ivl_18644 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3856
  signal tmp_ivl_18649 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3856
  signal tmp_ivl_1865 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3004
  signal tmp_ivl_18652 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3856
  signal tmp_ivl_18654 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3856
  signal tmp_ivl_18655 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3856
  signal tmp_ivl_18660 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3856
  signal tmp_ivl_18662 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3856
  signal tmp_ivl_18668 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3857
  signal tmp_ivl_18669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3857
  signal tmp_ivl_18674 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3857
  signal tmp_ivl_18677 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3857
  signal tmp_ivl_18679 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3857
  signal tmp_ivl_1868 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3004
  signal tmp_ivl_18680 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3857
  signal tmp_ivl_18685 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3857
  signal tmp_ivl_18687 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3857
  signal tmp_ivl_18693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3858
  signal tmp_ivl_18695 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3858
  signal tmp_ivl_18696 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3858
  signal tmp_ivl_1870 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3004
  signal tmp_ivl_18701 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3858
  signal tmp_ivl_18703 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3858
  signal tmp_ivl_18708 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3858
  signal tmp_ivl_1871 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3004
  signal tmp_ivl_18710 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3858
  signal tmp_ivl_18715 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3859
  signal tmp_ivl_18720 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3859
  signal tmp_ivl_18722 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3859
  signal tmp_ivl_18727 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3859
  signal tmp_ivl_18729 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3859
  signal tmp_ivl_18734 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3860
  signal tmp_ivl_18739 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3860
  signal tmp_ivl_18741 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3860
  signal tmp_ivl_18746 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3860
  signal tmp_ivl_18748 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3860
  signal tmp_ivl_18750 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3860
  signal tmp_ivl_18752 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3860
  signal tmp_ivl_18757 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3861
  signal tmp_ivl_1876 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3004
  signal tmp_ivl_18762 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3861
  signal tmp_ivl_18764 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3861
  signal tmp_ivl_18769 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3861
  signal tmp_ivl_18771 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3861
  signal tmp_ivl_18776 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3862
  signal tmp_ivl_1878 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3004
  signal tmp_ivl_18781 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3862
  signal tmp_ivl_18783 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3862
  signal tmp_ivl_18788 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3862
  signal tmp_ivl_18790 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3862
  signal tmp_ivl_18795 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3863
  signal tmp_ivl_188 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2946
  signal tmp_ivl_1880 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3004
  signal tmp_ivl_18800 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3863
  signal tmp_ivl_18802 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3863
  signal tmp_ivl_18807 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3863
  signal tmp_ivl_18809 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3863
  signal tmp_ivl_18815 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3864
  signal tmp_ivl_18816 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3864
  signal tmp_ivl_18821 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3864
  signal tmp_ivl_18824 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3864
  signal tmp_ivl_18826 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3864
  signal tmp_ivl_18827 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3864
  signal tmp_ivl_18832 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3864
  signal tmp_ivl_18834 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3864
  signal tmp_ivl_18839 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3865
  signal tmp_ivl_18844 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3865
  signal tmp_ivl_18846 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3865
  signal tmp_ivl_18851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3865
  signal tmp_ivl_18853 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3865
  signal tmp_ivl_18858 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3866
  signal tmp_ivl_1886 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3005
  signal tmp_ivl_18863 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3866
  signal tmp_ivl_18865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3866
  signal tmp_ivl_18870 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3866
  signal tmp_ivl_18872 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3866
  signal tmp_ivl_18874 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3866
  signal tmp_ivl_18876 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3866
  signal tmp_ivl_1888 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3005
  signal tmp_ivl_18881 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3867
  signal tmp_ivl_18886 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3867
  signal tmp_ivl_18888 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3867
  signal tmp_ivl_1889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3005
  signal tmp_ivl_18893 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3867
  signal tmp_ivl_18895 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3867
  signal tmp_ivl_189 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2946
  signal tmp_ivl_18901 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3868
  signal tmp_ivl_18902 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3868
  signal tmp_ivl_18907 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3868
  signal tmp_ivl_18910 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3868
  signal tmp_ivl_18912 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3868
  signal tmp_ivl_18913 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3868
  signal tmp_ivl_18918 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3868
  signal tmp_ivl_18920 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3868
  signal tmp_ivl_18926 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3869
  signal tmp_ivl_18928 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3869
  signal tmp_ivl_18929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3869
  signal tmp_ivl_18934 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3869
  signal tmp_ivl_18936 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3869
  signal tmp_ivl_1894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3005
  signal tmp_ivl_18941 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3869
  signal tmp_ivl_18943 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3869
  signal tmp_ivl_18948 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3870
  signal tmp_ivl_18953 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3870
  signal tmp_ivl_18955 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3870
  signal tmp_ivl_18960 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3870
  signal tmp_ivl_18962 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3870
  signal tmp_ivl_18967 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3871
  signal tmp_ivl_1897 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3005
  signal tmp_ivl_18972 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3871
  signal tmp_ivl_18974 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3871
  signal tmp_ivl_18979 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3871
  signal tmp_ivl_18981 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3871
  signal tmp_ivl_18983 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3871
  signal tmp_ivl_18985 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3871
  signal tmp_ivl_1899 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3005
  signal tmp_ivl_18990 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3872
  signal tmp_ivl_18995 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3872
  signal tmp_ivl_18997 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3872
  signal tmp_ivl_1900 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3005
  signal tmp_ivl_19002 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3872
  signal tmp_ivl_19004 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3872
  signal tmp_ivl_19010 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3873
  signal tmp_ivl_19011 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3873
  signal tmp_ivl_19016 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3873
  signal tmp_ivl_19019 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3873
  signal tmp_ivl_19021 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3873
  signal tmp_ivl_19022 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3873
  signal tmp_ivl_19027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3873
  signal tmp_ivl_19029 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3873
  signal tmp_ivl_19035 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3874
  signal tmp_ivl_19037 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3874
  signal tmp_ivl_19038 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3874
  signal tmp_ivl_19043 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3874
  signal tmp_ivl_19045 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3874
  signal tmp_ivl_1905 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3005
  signal tmp_ivl_19050 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3874
  signal tmp_ivl_19052 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3874
  signal tmp_ivl_19057 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3875
  signal tmp_ivl_19062 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3875
  signal tmp_ivl_19064 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3875
  signal tmp_ivl_19069 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3875
  signal tmp_ivl_1907 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3005
  signal tmp_ivl_19071 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3875
  signal tmp_ivl_19076 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3876
  signal tmp_ivl_19081 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3876
  signal tmp_ivl_19083 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3876
  signal tmp_ivl_19088 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3876
  signal tmp_ivl_1909 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3005
  signal tmp_ivl_19090 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3876
  signal tmp_ivl_19092 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3876
  signal tmp_ivl_19094 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3876
  signal tmp_ivl_19100 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3877
  signal tmp_ivl_19102 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3877
  signal tmp_ivl_19103 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3877
  signal tmp_ivl_19108 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3877
  signal tmp_ivl_19111 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3877
  signal tmp_ivl_19112 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3877
  signal tmp_ivl_19117 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3877
  signal tmp_ivl_19119 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3877
  signal tmp_ivl_19124 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3878
  signal tmp_ivl_19129 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3878
  signal tmp_ivl_19131 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3878
  signal tmp_ivl_19136 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3878
  signal tmp_ivl_19138 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3878
  signal tmp_ivl_19143 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3879
  signal tmp_ivl_19148 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3879
  signal tmp_ivl_1915 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3006
  signal tmp_ivl_19150 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3879
  signal tmp_ivl_19155 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3879
  signal tmp_ivl_19157 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3879
  signal tmp_ivl_19162 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3880
  signal tmp_ivl_19167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3880
  signal tmp_ivl_19169 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3880
  signal tmp_ivl_1917 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3006
  signal tmp_ivl_19174 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3880
  signal tmp_ivl_19176 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3880
  signal tmp_ivl_1918 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3006
  signal tmp_ivl_19181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3881
  signal tmp_ivl_19186 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3881
  signal tmp_ivl_19188 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3881
  signal tmp_ivl_19193 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3881
  signal tmp_ivl_19195 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3881
  signal tmp_ivl_19200 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3882
  signal tmp_ivl_19205 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3882
  signal tmp_ivl_19207 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3882
  signal tmp_ivl_19212 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3882
  signal tmp_ivl_19214 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3882
  signal tmp_ivl_19216 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3882
  signal tmp_ivl_19218 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3882
  signal tmp_ivl_19223 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3883
  signal tmp_ivl_19228 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3883
  signal tmp_ivl_1923 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3006
  signal tmp_ivl_19230 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3883
  signal tmp_ivl_19235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3883
  signal tmp_ivl_19237 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3883
  signal tmp_ivl_19243 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3884
  signal tmp_ivl_19245 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3884
  signal tmp_ivl_19246 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3884
  signal tmp_ivl_19251 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3884
  signal tmp_ivl_19253 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3884
  signal tmp_ivl_19258 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3884
  signal tmp_ivl_1926 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3006
  signal tmp_ivl_19260 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3884
  signal tmp_ivl_19265 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3885
  signal tmp_ivl_19270 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3885
  signal tmp_ivl_19272 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3885
  signal tmp_ivl_19277 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3885
  signal tmp_ivl_19279 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3885
  signal tmp_ivl_1928 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3006
  signal tmp_ivl_19281 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3885
  signal tmp_ivl_19283 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3885
  signal tmp_ivl_19288 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3886
  signal tmp_ivl_1929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3006
  signal tmp_ivl_19293 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3886
  signal tmp_ivl_19295 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3886
  signal tmp_ivl_19300 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3886
  signal tmp_ivl_19302 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3886
  signal tmp_ivl_19307 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3887
  signal tmp_ivl_19312 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3887
  signal tmp_ivl_19314 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3887
  signal tmp_ivl_19319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3887
  signal tmp_ivl_19321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3887
  signal tmp_ivl_19327 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3888
  signal tmp_ivl_19328 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3888
  signal tmp_ivl_19333 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3888
  signal tmp_ivl_19336 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3888
  signal tmp_ivl_19338 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3888
  signal tmp_ivl_19339 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3888
  signal tmp_ivl_1934 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3006
  signal tmp_ivl_19344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3888
  signal tmp_ivl_19346 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3888
  signal tmp_ivl_19351 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3889
  signal tmp_ivl_19356 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3889
  signal tmp_ivl_19358 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3889
  signal tmp_ivl_1936 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3006
  signal tmp_ivl_19363 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3889
  signal tmp_ivl_19365 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3889
  signal tmp_ivl_19370 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3890
  signal tmp_ivl_19375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3890
  signal tmp_ivl_19377 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3890
  signal tmp_ivl_1938 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3006
  signal tmp_ivl_19382 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3890
  signal tmp_ivl_19384 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3890
  signal tmp_ivl_19386 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3890
  signal tmp_ivl_19388 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3890
  signal tmp_ivl_19393 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3891
  signal tmp_ivl_19398 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3891
  signal tmp_ivl_194 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2946
  signal tmp_ivl_19400 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3891
  signal tmp_ivl_19405 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3891
  signal tmp_ivl_19407 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3891
  signal tmp_ivl_19413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3892
  signal tmp_ivl_19414 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3892
  signal tmp_ivl_19419 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3892
  signal tmp_ivl_19421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3892
  signal tmp_ivl_19426 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3892
  signal tmp_ivl_19428 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3892
  signal tmp_ivl_19433 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3893
  signal tmp_ivl_19438 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3893
  signal tmp_ivl_1944 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3007
  signal tmp_ivl_19440 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3893
  signal tmp_ivl_19445 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3893
  signal tmp_ivl_19447 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3893
  signal tmp_ivl_19452 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3894
  signal tmp_ivl_19457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3894
  signal tmp_ivl_19459 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3894
  signal tmp_ivl_1946 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3007
  signal tmp_ivl_19464 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3894
  signal tmp_ivl_19466 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3894
  signal tmp_ivl_19468 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3894
  signal tmp_ivl_1947 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3007
  signal tmp_ivl_19470 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3894
  signal tmp_ivl_19475 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3895
  signal tmp_ivl_19480 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3895
  signal tmp_ivl_19482 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3895
  signal tmp_ivl_19487 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3895
  signal tmp_ivl_19489 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3895
  signal tmp_ivl_19494 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3896
  signal tmp_ivl_19499 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3896
  signal tmp_ivl_19501 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3896
  signal tmp_ivl_19506 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3896
  signal tmp_ivl_19508 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3896
  signal tmp_ivl_19514 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3897
  signal tmp_ivl_19515 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3897
  signal tmp_ivl_1952 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3007
  signal tmp_ivl_19520 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3897
  signal tmp_ivl_19523 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3897
  signal tmp_ivl_19525 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3897
  signal tmp_ivl_19526 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3897
  signal tmp_ivl_19531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3897
  signal tmp_ivl_19533 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3897
  signal tmp_ivl_19538 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3898
  signal tmp_ivl_19543 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3898
  signal tmp_ivl_19545 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3898
  signal tmp_ivl_1955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3007
  signal tmp_ivl_19550 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3898
  signal tmp_ivl_19552 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3898
  signal tmp_ivl_19557 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3899
  signal tmp_ivl_19562 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3899
  signal tmp_ivl_19564 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3899
  signal tmp_ivl_19569 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3899
  signal tmp_ivl_1957 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3007
  signal tmp_ivl_19571 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3899
  signal tmp_ivl_19573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3899
  signal tmp_ivl_19575 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3899
  signal tmp_ivl_1958 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3007
  signal tmp_ivl_19580 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3900
  signal tmp_ivl_19585 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3900
  signal tmp_ivl_19587 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3900
  signal tmp_ivl_19592 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3900
  signal tmp_ivl_19594 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3900
  signal tmp_ivl_196 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2946
  signal tmp_ivl_19600 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3901
  signal tmp_ivl_19601 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3901
  signal tmp_ivl_19606 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3901
  signal tmp_ivl_19609 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3901
  signal tmp_ivl_19611 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3901
  signal tmp_ivl_19612 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3901
  signal tmp_ivl_19617 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3901
  signal tmp_ivl_19619 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3901
  signal tmp_ivl_19625 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3902
  signal tmp_ivl_19627 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3902
  signal tmp_ivl_19628 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3902
  signal tmp_ivl_1963 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3007
  signal tmp_ivl_19633 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3902
  signal tmp_ivl_19635 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3902
  signal tmp_ivl_19640 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3902
  signal tmp_ivl_19642 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3902
  signal tmp_ivl_19647 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3903
  signal tmp_ivl_1965 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3007
  signal tmp_ivl_19652 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3903
  signal tmp_ivl_19654 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3903
  signal tmp_ivl_19659 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3903
  signal tmp_ivl_19661 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3903
  signal tmp_ivl_19666 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3904
  signal tmp_ivl_1967 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3007
  signal tmp_ivl_19671 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3904
  signal tmp_ivl_19673 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3904
  signal tmp_ivl_19678 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3904
  signal tmp_ivl_19680 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3904
  signal tmp_ivl_19682 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3904
  signal tmp_ivl_19684 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3904
  signal tmp_ivl_19689 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3905
  signal tmp_ivl_19694 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3905
  signal tmp_ivl_19696 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3905
  signal tmp_ivl_19701 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3905
  signal tmp_ivl_19703 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3905
  signal tmp_ivl_19709 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3906
  signal tmp_ivl_19711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3906
  signal tmp_ivl_19712 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3906
  signal tmp_ivl_19717 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3906
  signal tmp_ivl_19720 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3906
  signal tmp_ivl_19721 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3906
  signal tmp_ivl_19726 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3906
  signal tmp_ivl_19728 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3906
  signal tmp_ivl_1973 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3008
  signal tmp_ivl_19733 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3907
  signal tmp_ivl_19738 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3907
  signal tmp_ivl_19740 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3907
  signal tmp_ivl_19745 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3907
  signal tmp_ivl_19747 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3907
  signal tmp_ivl_1975 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3008
  signal tmp_ivl_19752 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3908
  signal tmp_ivl_19757 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3908
  signal tmp_ivl_19759 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3908
  signal tmp_ivl_1976 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3008
  signal tmp_ivl_19764 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3908
  signal tmp_ivl_19766 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3908
  signal tmp_ivl_19768 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3908
  signal tmp_ivl_19770 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3908
  signal tmp_ivl_19775 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3909
  signal tmp_ivl_19780 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3909
  signal tmp_ivl_19782 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3909
  signal tmp_ivl_19787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3909
  signal tmp_ivl_19789 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3909
  signal tmp_ivl_19795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3910
  signal tmp_ivl_19797 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3910
  signal tmp_ivl_19798 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3910
  signal tmp_ivl_198 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2946
  signal tmp_ivl_19803 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3910
  signal tmp_ivl_19805 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3910
  signal tmp_ivl_1981 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3008
  signal tmp_ivl_19810 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3910
  signal tmp_ivl_19812 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3910
  signal tmp_ivl_19817 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3911
  signal tmp_ivl_19822 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3911
  signal tmp_ivl_19824 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3911
  signal tmp_ivl_19829 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3911
  signal tmp_ivl_19831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3911
  signal tmp_ivl_19833 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3911
  signal tmp_ivl_19835 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3911
  signal tmp_ivl_1984 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3008
  signal tmp_ivl_19840 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3912
  signal tmp_ivl_19845 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3912
  signal tmp_ivl_19847 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3912
  signal tmp_ivl_19852 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3912
  signal tmp_ivl_19854 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3912
  signal tmp_ivl_19859 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3913
  signal tmp_ivl_1986 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3008
  signal tmp_ivl_19864 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3913
  signal tmp_ivl_19866 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3913
  signal tmp_ivl_1987 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3008
  signal tmp_ivl_19871 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3913
  signal tmp_ivl_19873 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3913
  signal tmp_ivl_19875 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3913
  signal tmp_ivl_19877 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3913
  signal tmp_ivl_19882 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3914
  signal tmp_ivl_19887 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3914
  signal tmp_ivl_19889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3914
  signal tmp_ivl_19894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3914
  signal tmp_ivl_19896 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3914
  signal tmp_ivl_19901 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3915
  signal tmp_ivl_19906 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3915
  signal tmp_ivl_19908 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3915
  signal tmp_ivl_19913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3915
  signal tmp_ivl_19915 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3915
  signal tmp_ivl_19917 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3915
  signal tmp_ivl_19919 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3915
  signal tmp_ivl_1992 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3008
  signal tmp_ivl_19924 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3916
  signal tmp_ivl_19929 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3916
  signal tmp_ivl_19931 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3916
  signal tmp_ivl_19936 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3916
  signal tmp_ivl_19938 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3916
  signal tmp_ivl_1994 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3008
  signal tmp_ivl_19944 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3917
  signal tmp_ivl_19945 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3917
  signal tmp_ivl_19950 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3917
  signal tmp_ivl_19953 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3917
  signal tmp_ivl_19955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3917
  signal tmp_ivl_19956 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3917
  signal tmp_ivl_1996 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3008
  signal tmp_ivl_19961 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3917
  signal tmp_ivl_19963 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3917
  signal tmp_ivl_19968 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3918
  signal tmp_ivl_19973 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3918
  signal tmp_ivl_19975 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3918
  signal tmp_ivl_19980 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3918
  signal tmp_ivl_19982 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3918
  signal tmp_ivl_19987 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3919
  signal tmp_ivl_19992 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3919
  signal tmp_ivl_19994 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3919
  signal tmp_ivl_19999 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3919
  signal tmp_ivl_20 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2940
  signal tmp_ivl_20001 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3919
  signal tmp_ivl_20003 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3919
  signal tmp_ivl_20005 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3919
  signal tmp_ivl_20010 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3920
  signal tmp_ivl_20015 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3920
  signal tmp_ivl_20017 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3920
  signal tmp_ivl_2002 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3009
  signal tmp_ivl_20022 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3920
  signal tmp_ivl_20024 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3920
  signal tmp_ivl_20029 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3921
  signal tmp_ivl_20034 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3921
  signal tmp_ivl_20036 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3921
  signal tmp_ivl_2004 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3009
  signal tmp_ivl_20041 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3921
  signal tmp_ivl_20043 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3921
  signal tmp_ivl_20045 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3921
  signal tmp_ivl_20047 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3921
  signal tmp_ivl_2005 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3009
  signal tmp_ivl_20052 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3922
  signal tmp_ivl_20057 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3922
  signal tmp_ivl_20059 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3922
  signal tmp_ivl_20064 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3922
  signal tmp_ivl_20066 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3922
  signal tmp_ivl_20072 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3923
  signal tmp_ivl_20073 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3923
  signal tmp_ivl_20078 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3923
  signal tmp_ivl_20081 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3923
  signal tmp_ivl_20083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3923
  signal tmp_ivl_20084 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3923
  signal tmp_ivl_20089 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3923
  signal tmp_ivl_20091 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3923
  signal tmp_ivl_20097 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3924
  signal tmp_ivl_20099 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3924
  signal tmp_ivl_2010 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3009
  signal tmp_ivl_20100 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3924
  signal tmp_ivl_20105 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3924
  signal tmp_ivl_20107 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3924
  signal tmp_ivl_20112 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3924
  signal tmp_ivl_20114 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3924
  signal tmp_ivl_20119 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3925
  signal tmp_ivl_20124 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3925
  signal tmp_ivl_20126 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3925
  signal tmp_ivl_2013 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3009
  signal tmp_ivl_20131 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3925
  signal tmp_ivl_20133 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3925
  signal tmp_ivl_20138 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3926
  signal tmp_ivl_20143 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3926
  signal tmp_ivl_20145 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3926
  signal tmp_ivl_2015 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3009
  signal tmp_ivl_20150 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3926
  signal tmp_ivl_20152 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3926
  signal tmp_ivl_20154 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3926
  signal tmp_ivl_20156 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3926
  signal tmp_ivl_2016 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3009
  signal tmp_ivl_20161 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3927
  signal tmp_ivl_20166 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3927
  signal tmp_ivl_20168 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3927
  signal tmp_ivl_20173 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3927
  signal tmp_ivl_20175 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3927
  signal tmp_ivl_20180 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3928
  signal tmp_ivl_20185 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3928
  signal tmp_ivl_20187 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3928
  signal tmp_ivl_20192 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3928
  signal tmp_ivl_20194 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3928
  signal tmp_ivl_20196 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3928
  signal tmp_ivl_20198 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3928
  signal tmp_ivl_20203 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3929
  signal tmp_ivl_20208 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3929
  signal tmp_ivl_2021 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3009
  signal tmp_ivl_20210 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3929
  signal tmp_ivl_20215 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3929
  signal tmp_ivl_20217 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3929
  signal tmp_ivl_20223 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3930
  signal tmp_ivl_20224 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3930
  signal tmp_ivl_20229 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3930
  signal tmp_ivl_2023 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3009
  signal tmp_ivl_20232 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3930
  signal tmp_ivl_20234 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3930
  signal tmp_ivl_20235 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3930
  signal tmp_ivl_20240 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3930
  signal tmp_ivl_20242 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3930
  signal tmp_ivl_20247 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3931
  signal tmp_ivl_2025 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3009
  signal tmp_ivl_20252 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3931
  signal tmp_ivl_20254 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3931
  signal tmp_ivl_20259 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3931
  signal tmp_ivl_20261 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3931
  signal tmp_ivl_20266 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3932
  signal tmp_ivl_20271 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3932
  signal tmp_ivl_20273 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3932
  signal tmp_ivl_20278 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3932
  signal tmp_ivl_20280 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3932
  signal tmp_ivl_20282 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3932
  signal tmp_ivl_20284 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3932
  signal tmp_ivl_20289 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3933
  signal tmp_ivl_20294 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3933
  signal tmp_ivl_20296 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3933
  signal tmp_ivl_20301 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3933
  signal tmp_ivl_20303 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3933
  signal tmp_ivl_20309 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3934
  signal tmp_ivl_2031 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3010
  signal tmp_ivl_20310 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3934
  signal tmp_ivl_20315 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3934
  signal tmp_ivl_20318 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3934
  signal tmp_ivl_20320 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3934
  signal tmp_ivl_20321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3934
  signal tmp_ivl_20326 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3934
  signal tmp_ivl_20328 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3934
  signal tmp_ivl_2033 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3010
  signal tmp_ivl_20334 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3935
  signal tmp_ivl_20336 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3935
  signal tmp_ivl_20337 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3935
  signal tmp_ivl_2034 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3010
  signal tmp_ivl_20342 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3935
  signal tmp_ivl_20344 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3935
  signal tmp_ivl_20349 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3935
  signal tmp_ivl_20351 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3935
  signal tmp_ivl_20356 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3936
  signal tmp_ivl_20361 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3936
  signal tmp_ivl_20363 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3936
  signal tmp_ivl_20368 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3936
  signal tmp_ivl_20370 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3936
  signal tmp_ivl_20375 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3937
  signal tmp_ivl_20380 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3937
  signal tmp_ivl_20382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3937
  signal tmp_ivl_20387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3937
  signal tmp_ivl_20389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3937
  signal tmp_ivl_2039 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3010
  signal tmp_ivl_20391 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3937
  signal tmp_ivl_20393 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3937
  signal tmp_ivl_20398 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3938
  signal tmp_ivl_204 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2947
  signal tmp_ivl_20403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3938
  signal tmp_ivl_20405 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3938
  signal tmp_ivl_20410 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3938
  signal tmp_ivl_20412 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3938
  signal tmp_ivl_20418 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3939
  signal tmp_ivl_2042 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3010
  signal tmp_ivl_20420 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3939
  signal tmp_ivl_20421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3939
  signal tmp_ivl_20426 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3939
  signal tmp_ivl_20429 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3939
  signal tmp_ivl_20430 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3939
  signal tmp_ivl_20435 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3939
  signal tmp_ivl_20437 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3939
  signal tmp_ivl_2044 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3010
  signal tmp_ivl_20442 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3940
  signal tmp_ivl_20447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3940
  signal tmp_ivl_20449 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3940
  signal tmp_ivl_2045 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3010
  signal tmp_ivl_20454 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3940
  signal tmp_ivl_20456 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3940
  signal tmp_ivl_20461 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3941
  signal tmp_ivl_20466 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3941
  signal tmp_ivl_20468 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3941
  signal tmp_ivl_20473 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3941
  signal tmp_ivl_20475 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3941
  signal tmp_ivl_20477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3941
  signal tmp_ivl_20479 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3941
  signal tmp_ivl_20484 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3942
  signal tmp_ivl_20489 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3942
  signal tmp_ivl_20491 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3942
  signal tmp_ivl_20496 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3942
  signal tmp_ivl_20498 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3942
  signal tmp_ivl_2050 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3010
  signal tmp_ivl_20503 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3943
  signal tmp_ivl_20508 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3943
  signal tmp_ivl_20510 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3943
  signal tmp_ivl_20515 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3943
  signal tmp_ivl_20517 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3943
  signal tmp_ivl_20519 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3943
  signal tmp_ivl_2052 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3010
  signal tmp_ivl_20521 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3943
  signal tmp_ivl_20526 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3944
  signal tmp_ivl_20531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3944
  signal tmp_ivl_20533 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3944
  signal tmp_ivl_20538 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3944
  signal tmp_ivl_2054 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3010
  signal tmp_ivl_20540 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3944
  signal tmp_ivl_20546 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3945
  signal tmp_ivl_20548 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3945
  signal tmp_ivl_20549 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3945
  signal tmp_ivl_20554 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3945
  signal tmp_ivl_20556 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3945
  signal tmp_ivl_20561 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3945
  signal tmp_ivl_20563 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3945
  signal tmp_ivl_20568 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3946
  signal tmp_ivl_20573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3946
  signal tmp_ivl_20575 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3946
  signal tmp_ivl_20580 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3946
  signal tmp_ivl_20582 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3946
  signal tmp_ivl_20584 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3946
  signal tmp_ivl_20586 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3946
  signal tmp_ivl_20591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3947
  signal tmp_ivl_20596 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3947
  signal tmp_ivl_20598 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3947
  signal tmp_ivl_206 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2947
  signal tmp_ivl_2060 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3011
  signal tmp_ivl_20603 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3947
  signal tmp_ivl_20605 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3947
  signal tmp_ivl_20610 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3948
  signal tmp_ivl_20615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3948
  signal tmp_ivl_20617 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3948
  signal tmp_ivl_2062 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3011
  signal tmp_ivl_20622 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3948
  signal tmp_ivl_20624 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3948
  signal tmp_ivl_20626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3948
  signal tmp_ivl_20628 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3948
  signal tmp_ivl_2063 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3011
  signal tmp_ivl_20633 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3949
  signal tmp_ivl_20638 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3949
  signal tmp_ivl_20640 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3949
  signal tmp_ivl_20645 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3949
  signal tmp_ivl_20647 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3949
  signal tmp_ivl_20652 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3950
  signal tmp_ivl_20657 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3950
  signal tmp_ivl_20659 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3950
  signal tmp_ivl_20664 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3950
  signal tmp_ivl_20666 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3950
  signal tmp_ivl_20668 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3950
  signal tmp_ivl_20670 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3950
  signal tmp_ivl_20675 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3951
  signal tmp_ivl_2068 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3011
  signal tmp_ivl_20680 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3951
  signal tmp_ivl_20682 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3951
  signal tmp_ivl_20687 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3951
  signal tmp_ivl_20689 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3951
  signal tmp_ivl_20695 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3952
  signal tmp_ivl_20696 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3952
  signal tmp_ivl_207 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2947
  signal tmp_ivl_20701 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3952
  signal tmp_ivl_20704 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3952
  signal tmp_ivl_20706 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3952
  signal tmp_ivl_20707 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3952
  signal tmp_ivl_2071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3011
  signal tmp_ivl_20712 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3952
  signal tmp_ivl_20714 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3952
  signal tmp_ivl_20719 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3953
  signal tmp_ivl_20724 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3953
  signal tmp_ivl_20726 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3953
  signal tmp_ivl_2073 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3011
  signal tmp_ivl_20731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3953
  signal tmp_ivl_20733 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3953
  signal tmp_ivl_20738 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3954
  signal tmp_ivl_2074 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3011
  signal tmp_ivl_20743 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3954
  signal tmp_ivl_20745 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3954
  signal tmp_ivl_20750 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3954
  signal tmp_ivl_20752 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3954
  signal tmp_ivl_20754 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3954
  signal tmp_ivl_20756 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3954
  signal tmp_ivl_20761 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3955
  signal tmp_ivl_20766 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3955
  signal tmp_ivl_20768 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3955
  signal tmp_ivl_20773 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3955
  signal tmp_ivl_20775 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3955
  signal tmp_ivl_20780 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3956
  signal tmp_ivl_20785 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3956
  signal tmp_ivl_20787 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3956
  signal tmp_ivl_2079 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3011
  signal tmp_ivl_20792 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3956
  signal tmp_ivl_20794 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3956
  signal tmp_ivl_20796 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3956
  signal tmp_ivl_20798 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3956
  signal tmp_ivl_20803 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3957
  signal tmp_ivl_20808 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3957
  signal tmp_ivl_2081 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3011
  signal tmp_ivl_20810 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3957
  signal tmp_ivl_20815 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3957
  signal tmp_ivl_20817 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3957
  signal tmp_ivl_20823 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3958
  signal tmp_ivl_20824 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3958
  signal tmp_ivl_20829 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3958
  signal tmp_ivl_2083 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3011
  signal tmp_ivl_20832 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3958
  signal tmp_ivl_20834 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3958
  signal tmp_ivl_20835 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3958
  signal tmp_ivl_20840 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3958
  signal tmp_ivl_20842 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3958
  signal tmp_ivl_20848 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3959
  signal tmp_ivl_20850 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3959
  signal tmp_ivl_20851 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3959
  signal tmp_ivl_20856 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3959
  signal tmp_ivl_20858 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3959
  signal tmp_ivl_20863 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3959
  signal tmp_ivl_20865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3959
  signal tmp_ivl_20870 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3960
  signal tmp_ivl_20875 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3960
  signal tmp_ivl_20877 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3960
  signal tmp_ivl_20882 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3960
  signal tmp_ivl_20884 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3960
  signal tmp_ivl_20889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3961
  signal tmp_ivl_2089 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3012
  signal tmp_ivl_20894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3961
  signal tmp_ivl_20896 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3961
  signal tmp_ivl_20901 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3961
  signal tmp_ivl_20903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3961
  signal tmp_ivl_20905 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3961
  signal tmp_ivl_20907 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3961
  signal tmp_ivl_2091 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3012
  signal tmp_ivl_20912 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3962
  signal tmp_ivl_20917 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3962
  signal tmp_ivl_20919 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3962
  signal tmp_ivl_2092 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3012
  signal tmp_ivl_20924 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3962
  signal tmp_ivl_20926 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3962
  signal tmp_ivl_20931 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3963
  signal tmp_ivl_20936 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3963
  signal tmp_ivl_20938 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3963
  signal tmp_ivl_20943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3963
  signal tmp_ivl_20945 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3963
  signal tmp_ivl_20947 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3963
  signal tmp_ivl_20949 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3963
  signal tmp_ivl_20954 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3964
  signal tmp_ivl_20959 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3964
  signal tmp_ivl_20961 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3964
  signal tmp_ivl_20966 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3964
  signal tmp_ivl_20968 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3964
  signal tmp_ivl_2097 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3012
  signal tmp_ivl_20974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3965
  signal tmp_ivl_20976 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3965
  signal tmp_ivl_20977 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3965
  signal tmp_ivl_20982 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3965
  signal tmp_ivl_20985 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3965
  signal tmp_ivl_20986 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3965
  signal tmp_ivl_20991 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3965
  signal tmp_ivl_20993 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3965
  signal tmp_ivl_20998 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3966
  signal tmp_ivl_2100 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3012
  signal tmp_ivl_21003 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3966
  signal tmp_ivl_21005 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3966
  signal tmp_ivl_21010 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3966
  signal tmp_ivl_21012 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3966
  signal tmp_ivl_21017 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3967
  signal tmp_ivl_2102 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3012
  signal tmp_ivl_21022 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3967
  signal tmp_ivl_21024 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3967
  signal tmp_ivl_21029 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3967
  signal tmp_ivl_2103 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3012
  signal tmp_ivl_21031 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3967
  signal tmp_ivl_21036 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3968
  signal tmp_ivl_21041 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3968
  signal tmp_ivl_21043 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3968
  signal tmp_ivl_21048 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3968
  signal tmp_ivl_21050 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3968
  signal tmp_ivl_21055 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3969
  signal tmp_ivl_21060 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3969
  signal tmp_ivl_21062 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3969
  signal tmp_ivl_21067 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3969
  signal tmp_ivl_21069 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3969
  signal tmp_ivl_21071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3969
  signal tmp_ivl_21073 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3969
  signal tmp_ivl_21078 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3970
  signal tmp_ivl_2108 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3012
  signal tmp_ivl_21083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3970
  signal tmp_ivl_21085 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3970
  signal tmp_ivl_21090 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3970
  signal tmp_ivl_21092 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3970
  signal tmp_ivl_21098 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3971
  signal tmp_ivl_2110 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3012
  signal tmp_ivl_21100 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3971
  signal tmp_ivl_21101 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3971
  signal tmp_ivl_21106 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3971
  signal tmp_ivl_21108 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3971
  signal tmp_ivl_21113 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3971
  signal tmp_ivl_21115 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3971
  signal tmp_ivl_2112 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3012
  signal tmp_ivl_21120 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3972
  signal tmp_ivl_21125 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3972
  signal tmp_ivl_21127 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3972
  signal tmp_ivl_21132 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3972
  signal tmp_ivl_21134 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3972
  signal tmp_ivl_21136 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3972
  signal tmp_ivl_21138 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3972
  signal tmp_ivl_21143 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3973
  signal tmp_ivl_21148 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3973
  signal tmp_ivl_21150 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3973
  signal tmp_ivl_21155 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3973
  signal tmp_ivl_21157 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3973
  signal tmp_ivl_21162 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3974
  signal tmp_ivl_21167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3974
  signal tmp_ivl_21169 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3974
  signal tmp_ivl_21174 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3974
  signal tmp_ivl_21176 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3974
  signal tmp_ivl_21178 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3974
  signal tmp_ivl_2118 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3013
  signal tmp_ivl_21180 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3974
  signal tmp_ivl_21185 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3975
  signal tmp_ivl_21190 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3975
  signal tmp_ivl_21192 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3975
  signal tmp_ivl_21197 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3975
  signal tmp_ivl_21199 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3975
  signal tmp_ivl_212 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2947
  signal tmp_ivl_2120 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3013
  signal tmp_ivl_21205 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3976
  signal tmp_ivl_21206 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3976
  signal tmp_ivl_2121 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3013
  signal tmp_ivl_21211 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3976
  signal tmp_ivl_21214 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3976
  signal tmp_ivl_21216 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3976
  signal tmp_ivl_21217 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3976
  signal tmp_ivl_21222 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3976
  signal tmp_ivl_21224 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3976
  signal tmp_ivl_21229 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3977
  signal tmp_ivl_21234 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3977
  signal tmp_ivl_21236 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3977
  signal tmp_ivl_21241 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3977
  signal tmp_ivl_21243 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3977
  signal tmp_ivl_21248 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3978
  signal tmp_ivl_21253 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3978
  signal tmp_ivl_21255 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3978
  signal tmp_ivl_2126 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3013
  signal tmp_ivl_21260 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3978
  signal tmp_ivl_21262 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3978
  signal tmp_ivl_21264 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3978
  signal tmp_ivl_21266 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3978
  signal tmp_ivl_21271 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3979
  signal tmp_ivl_21276 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3979
  signal tmp_ivl_21278 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3979
  signal tmp_ivl_21283 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3979
  signal tmp_ivl_21285 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3979
  signal tmp_ivl_2129 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3013
  signal tmp_ivl_21290 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3980
  signal tmp_ivl_21295 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3980
  signal tmp_ivl_21297 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3980
  signal tmp_ivl_21302 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3980
  signal tmp_ivl_21304 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3980
  signal tmp_ivl_21306 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3980
  signal tmp_ivl_21308 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3980
  signal tmp_ivl_2131 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3013
  signal tmp_ivl_21313 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3981
  signal tmp_ivl_21318 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3981
  signal tmp_ivl_2132 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3013
  signal tmp_ivl_21320 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3981
  signal tmp_ivl_21325 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3981
  signal tmp_ivl_21327 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3981
  signal tmp_ivl_21332 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3982
  signal tmp_ivl_21337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3982
  signal tmp_ivl_21339 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3982
  signal tmp_ivl_21344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3982
  signal tmp_ivl_21346 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3982
  signal tmp_ivl_21348 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3982
  signal tmp_ivl_21350 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3982
  signal tmp_ivl_21355 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3983
  signal tmp_ivl_21360 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3983
  signal tmp_ivl_21362 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3983
  signal tmp_ivl_21367 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3983
  signal tmp_ivl_21369 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3983
  signal tmp_ivl_2137 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3013
  signal tmp_ivl_21375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3984
  signal tmp_ivl_21376 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3984
  signal tmp_ivl_21381 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3984
  signal tmp_ivl_21383 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3984
  signal tmp_ivl_21388 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3984
  signal tmp_ivl_2139 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3013
  signal tmp_ivl_21390 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3984
  signal tmp_ivl_21395 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3985
  signal tmp_ivl_21400 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3985
  signal tmp_ivl_21402 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3985
  signal tmp_ivl_21407 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3985
  signal tmp_ivl_21409 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3985
  signal tmp_ivl_2141 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3013
  signal tmp_ivl_21414 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3986
  signal tmp_ivl_21419 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3986
  signal tmp_ivl_21421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3986
  signal tmp_ivl_21426 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3986
  signal tmp_ivl_21428 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3986
  signal tmp_ivl_21430 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3986
  signal tmp_ivl_21432 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3986
  signal tmp_ivl_21437 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3987
  signal tmp_ivl_21442 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3987
  signal tmp_ivl_21444 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3987
  signal tmp_ivl_21449 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3987
  signal tmp_ivl_21451 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3987
  signal tmp_ivl_21456 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3988
  signal tmp_ivl_21461 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3988
  signal tmp_ivl_21463 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3988
  signal tmp_ivl_21468 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3988
  signal tmp_ivl_2147 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3014
  signal tmp_ivl_21470 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3988
  signal tmp_ivl_21472 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3988
  signal tmp_ivl_21474 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3988
  signal tmp_ivl_21479 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3989
  signal tmp_ivl_21484 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3989
  signal tmp_ivl_21486 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3989
  signal tmp_ivl_2149 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3014
  signal tmp_ivl_21491 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3989
  signal tmp_ivl_21493 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3989
  signal tmp_ivl_21499 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3990
  signal tmp_ivl_215 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2947
  signal tmp_ivl_2150 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3014
  signal tmp_ivl_21500 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3990
  signal tmp_ivl_21505 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3990
  signal tmp_ivl_21508 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3990
  signal tmp_ivl_21510 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3990
  signal tmp_ivl_21511 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3990
  signal tmp_ivl_21516 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3990
  signal tmp_ivl_21518 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3990
  signal tmp_ivl_21523 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3991
  signal tmp_ivl_21528 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3991
  signal tmp_ivl_21530 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3991
  signal tmp_ivl_21535 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3991
  signal tmp_ivl_21537 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3991
  signal tmp_ivl_21542 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3992
  signal tmp_ivl_21547 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3992
  signal tmp_ivl_21549 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3992
  signal tmp_ivl_2155 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3014
  signal tmp_ivl_21554 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3992
  signal tmp_ivl_21556 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3992
  signal tmp_ivl_21558 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3992
  signal tmp_ivl_21560 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3992
  signal tmp_ivl_21565 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3993
  signal tmp_ivl_21570 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3993
  signal tmp_ivl_21572 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3993
  signal tmp_ivl_21577 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3993
  signal tmp_ivl_21579 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3993
  signal tmp_ivl_2158 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3014
  signal tmp_ivl_21584 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3994
  signal tmp_ivl_21589 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3994
  signal tmp_ivl_21591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3994
  signal tmp_ivl_21596 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3994
  signal tmp_ivl_21598 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3994
  signal tmp_ivl_2160 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3014
  signal tmp_ivl_21600 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3994
  signal tmp_ivl_21602 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3994
  signal tmp_ivl_21607 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3995
  signal tmp_ivl_2161 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3014
  signal tmp_ivl_21612 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3995
  signal tmp_ivl_21614 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3995
  signal tmp_ivl_21619 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3995
  signal tmp_ivl_21621 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3995
  signal tmp_ivl_21626 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3996
  signal tmp_ivl_21631 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3996
  signal tmp_ivl_21633 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3996
  signal tmp_ivl_21638 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3996
  signal tmp_ivl_21640 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3996
  signal tmp_ivl_21642 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3996
  signal tmp_ivl_21644 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3996
  signal tmp_ivl_21649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3997
  signal tmp_ivl_21654 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3997
  signal tmp_ivl_21656 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3997
  signal tmp_ivl_2166 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3014
  signal tmp_ivl_21661 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3997
  signal tmp_ivl_21663 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3997
  signal tmp_ivl_21669 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3998
  signal tmp_ivl_21670 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3998
  signal tmp_ivl_21675 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3998
  signal tmp_ivl_21678 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3998
  signal tmp_ivl_2168 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3014
  signal tmp_ivl_21680 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3998
  signal tmp_ivl_21681 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3998
  signal tmp_ivl_21686 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3998
  signal tmp_ivl_21688 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3998
  signal tmp_ivl_21694 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3999
  signal tmp_ivl_21696 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3999
  signal tmp_ivl_21697 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3999
  signal tmp_ivl_217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2947
  signal tmp_ivl_2170 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3014
  signal tmp_ivl_21702 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3999
  signal tmp_ivl_21704 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3999
  signal tmp_ivl_21709 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3999
  signal tmp_ivl_21711 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3999
  signal tmp_ivl_21716 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4000
  signal tmp_ivl_21721 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4000
  signal tmp_ivl_21723 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4000
  signal tmp_ivl_21728 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4000
  signal tmp_ivl_21730 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4000
  signal tmp_ivl_21735 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4001
  signal tmp_ivl_21740 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4001
  signal tmp_ivl_21742 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4001
  signal tmp_ivl_21747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4001
  signal tmp_ivl_21749 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4001
  signal tmp_ivl_21751 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4001
  signal tmp_ivl_21753 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4001
  signal tmp_ivl_21758 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4002
  signal tmp_ivl_2176 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3015
  signal tmp_ivl_21763 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4002
  signal tmp_ivl_21765 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4002
  signal tmp_ivl_21770 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4002
  signal tmp_ivl_21772 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4002
  signal tmp_ivl_21777 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4003
  signal tmp_ivl_2178 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3015
  signal tmp_ivl_21782 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4003
  signal tmp_ivl_21784 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4003
  signal tmp_ivl_21789 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4003
  signal tmp_ivl_2179 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3015
  signal tmp_ivl_21791 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4003
  signal tmp_ivl_21793 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4003
  signal tmp_ivl_21795 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4003
  signal tmp_ivl_218 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2947
  signal tmp_ivl_21800 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4004
  signal tmp_ivl_21805 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4004
  signal tmp_ivl_21807 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4004
  signal tmp_ivl_21812 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4004
  signal tmp_ivl_21814 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4004
  signal tmp_ivl_21820 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4005
  signal tmp_ivl_21822 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4005
  signal tmp_ivl_21823 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4005
  signal tmp_ivl_21828 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4005
  signal tmp_ivl_21831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4005
  signal tmp_ivl_21832 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4005
  signal tmp_ivl_21837 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4005
  signal tmp_ivl_21839 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4005
  signal tmp_ivl_2184 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3015
  signal tmp_ivl_21844 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4006
  signal tmp_ivl_21849 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4006
  signal tmp_ivl_21851 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4006
  signal tmp_ivl_21856 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4006
  signal tmp_ivl_21858 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4006
  signal tmp_ivl_21863 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4007
  signal tmp_ivl_21868 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4007
  signal tmp_ivl_2187 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3015
  signal tmp_ivl_21870 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4007
  signal tmp_ivl_21875 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4007
  signal tmp_ivl_21877 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4007
  signal tmp_ivl_21879 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4007
  signal tmp_ivl_21881 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4007
  signal tmp_ivl_21886 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4008
  signal tmp_ivl_2189 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3015
  signal tmp_ivl_21891 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4008
  signal tmp_ivl_21893 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4008
  signal tmp_ivl_21898 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4008
  signal tmp_ivl_2190 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3015
  signal tmp_ivl_21900 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4008
  signal tmp_ivl_21905 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4009
  signal tmp_ivl_21910 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4009
  signal tmp_ivl_21912 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4009
  signal tmp_ivl_21917 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4009
  signal tmp_ivl_21919 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4009
  signal tmp_ivl_21921 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4009
  signal tmp_ivl_21923 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4009
  signal tmp_ivl_21928 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4010
  signal tmp_ivl_21933 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4010
  signal tmp_ivl_21935 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4010
  signal tmp_ivl_21940 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4010
  signal tmp_ivl_21942 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4010
  signal tmp_ivl_21948 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4011
  signal tmp_ivl_2195 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3015
  signal tmp_ivl_21950 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4011
  signal tmp_ivl_21951 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4011
  signal tmp_ivl_21956 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4011
  signal tmp_ivl_21958 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4011
  signal tmp_ivl_21963 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4011
  signal tmp_ivl_21965 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4011
  signal tmp_ivl_2197 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3015
  signal tmp_ivl_21970 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4012
  signal tmp_ivl_21975 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4012
  signal tmp_ivl_21977 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4012
  signal tmp_ivl_21982 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4012
  signal tmp_ivl_21984 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4012
  signal tmp_ivl_21986 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4012
  signal tmp_ivl_21988 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4012
  signal tmp_ivl_2199 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3015
  signal tmp_ivl_21993 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4013
  signal tmp_ivl_21998 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4013
  signal tmp_ivl_22 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2940
  signal tmp_ivl_22000 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4013
  signal tmp_ivl_22005 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4013
  signal tmp_ivl_22007 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4013
  signal tmp_ivl_22012 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4014
  signal tmp_ivl_22017 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4014
  signal tmp_ivl_22019 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4014
  signal tmp_ivl_22024 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4014
  signal tmp_ivl_22026 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4014
  signal tmp_ivl_22028 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4014
  signal tmp_ivl_22030 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4014
  signal tmp_ivl_22035 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4015
  signal tmp_ivl_22040 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4015
  signal tmp_ivl_22042 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4015
  signal tmp_ivl_22047 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4015
  signal tmp_ivl_22049 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4015
  signal tmp_ivl_2205 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3016
  signal tmp_ivl_22054 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4016
  signal tmp_ivl_22059 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4016
  signal tmp_ivl_22061 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4016
  signal tmp_ivl_22066 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4016
  signal tmp_ivl_22068 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4016
  signal tmp_ivl_2207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3016
  signal tmp_ivl_22070 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4016
  signal tmp_ivl_22072 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4016
  signal tmp_ivl_22077 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4017
  signal tmp_ivl_2208 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3016
  signal tmp_ivl_22082 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4017
  signal tmp_ivl_22084 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4017
  signal tmp_ivl_22089 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4017
  signal tmp_ivl_22091 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4017
  signal tmp_ivl_22097 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4018
  signal tmp_ivl_22098 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4018
  signal tmp_ivl_22103 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4018
  signal tmp_ivl_22106 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4018
  signal tmp_ivl_22108 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4018
  signal tmp_ivl_22109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4018
  signal tmp_ivl_22114 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4018
  signal tmp_ivl_22116 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4018
  signal tmp_ivl_22121 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4019
  signal tmp_ivl_22126 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4019
  signal tmp_ivl_22128 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4019
  signal tmp_ivl_2213 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3016
  signal tmp_ivl_22133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4019
  signal tmp_ivl_22135 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4019
  signal tmp_ivl_22140 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4020
  signal tmp_ivl_22145 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4020
  signal tmp_ivl_22147 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4020
  signal tmp_ivl_22152 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4020
  signal tmp_ivl_22154 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4020
  signal tmp_ivl_22156 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4020
  signal tmp_ivl_22158 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4020
  signal tmp_ivl_2216 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3016
  signal tmp_ivl_22163 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4021
  signal tmp_ivl_22168 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4021
  signal tmp_ivl_22170 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4021
  signal tmp_ivl_22175 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4021
  signal tmp_ivl_22177 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4021
  signal tmp_ivl_2218 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3016
  signal tmp_ivl_22182 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4022
  signal tmp_ivl_22187 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4022
  signal tmp_ivl_22189 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4022
  signal tmp_ivl_2219 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3016
  signal tmp_ivl_22194 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4022
  signal tmp_ivl_22196 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4022
  signal tmp_ivl_22198 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4022
  signal tmp_ivl_22200 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4022
  signal tmp_ivl_22205 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4023
  signal tmp_ivl_22210 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4023
  signal tmp_ivl_22212 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4023
  signal tmp_ivl_22217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4023
  signal tmp_ivl_22219 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4023
  signal tmp_ivl_22224 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4024
  signal tmp_ivl_22229 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4024
  signal tmp_ivl_22231 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4024
  signal tmp_ivl_22236 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4024
  signal tmp_ivl_22238 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4024
  signal tmp_ivl_2224 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3016
  signal tmp_ivl_22240 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4024
  signal tmp_ivl_22242 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4024
  signal tmp_ivl_22247 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4025
  signal tmp_ivl_22252 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4025
  signal tmp_ivl_22254 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4025
  signal tmp_ivl_22259 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4025
  signal tmp_ivl_2226 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3016
  signal tmp_ivl_22261 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4025
  signal tmp_ivl_22267 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4026
  signal tmp_ivl_22268 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4026
  signal tmp_ivl_22273 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4026
  signal tmp_ivl_22276 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4026
  signal tmp_ivl_22278 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4026
  signal tmp_ivl_22279 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4026
  signal tmp_ivl_2228 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3016
  signal tmp_ivl_22284 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4026
  signal tmp_ivl_22286 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4026
  signal tmp_ivl_22292 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4027
  signal tmp_ivl_22294 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4027
  signal tmp_ivl_22295 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4027
  signal tmp_ivl_223 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2947
  signal tmp_ivl_22300 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4027
  signal tmp_ivl_22302 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4027
  signal tmp_ivl_22307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4027
  signal tmp_ivl_22309 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4027
  signal tmp_ivl_22314 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4028
  signal tmp_ivl_22319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4028
  signal tmp_ivl_22321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4028
  signal tmp_ivl_22326 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4028
  signal tmp_ivl_22328 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4028
  signal tmp_ivl_22333 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4029
  signal tmp_ivl_22338 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4029
  signal tmp_ivl_2234 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3017
  signal tmp_ivl_22340 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4029
  signal tmp_ivl_22345 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4029
  signal tmp_ivl_22347 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4029
  signal tmp_ivl_22349 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4029
  signal tmp_ivl_22351 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4029
  signal tmp_ivl_22356 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4030
  signal tmp_ivl_2236 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3017
  signal tmp_ivl_22361 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4030
  signal tmp_ivl_22363 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4030
  signal tmp_ivl_22368 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4030
  signal tmp_ivl_2237 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3017
  signal tmp_ivl_22370 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4030
  signal tmp_ivl_22375 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4031
  signal tmp_ivl_22380 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4031
  signal tmp_ivl_22382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4031
  signal tmp_ivl_22387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4031
  signal tmp_ivl_22389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4031
  signal tmp_ivl_22391 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4031
  signal tmp_ivl_22393 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4031
  signal tmp_ivl_22398 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4032
  signal tmp_ivl_22403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4032
  signal tmp_ivl_22405 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4032
  signal tmp_ivl_22410 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4032
  signal tmp_ivl_22412 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4032
  signal tmp_ivl_22417 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4033
  signal tmp_ivl_2242 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3017
  signal tmp_ivl_22422 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4033
  signal tmp_ivl_22424 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4033
  signal tmp_ivl_22429 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4033
  signal tmp_ivl_22431 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4033
  signal tmp_ivl_22433 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4033
  signal tmp_ivl_22435 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4033
  signal tmp_ivl_22440 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4034
  signal tmp_ivl_22445 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4034
  signal tmp_ivl_22447 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4034
  signal tmp_ivl_2245 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3017
  signal tmp_ivl_22452 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4034
  signal tmp_ivl_22454 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4034
  signal tmp_ivl_22460 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4035
  signal tmp_ivl_22461 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4035
  signal tmp_ivl_22466 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4035
  signal tmp_ivl_22469 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4035
  signal tmp_ivl_2247 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3017
  signal tmp_ivl_22471 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4035
  signal tmp_ivl_22472 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4035
  signal tmp_ivl_22477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4035
  signal tmp_ivl_22479 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4035
  signal tmp_ivl_2248 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3017
  signal tmp_ivl_22484 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4036
  signal tmp_ivl_22489 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4036
  signal tmp_ivl_22491 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4036
  signal tmp_ivl_22496 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4036
  signal tmp_ivl_22498 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4036
  signal tmp_ivl_225 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2947
  signal tmp_ivl_22503 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4037
  signal tmp_ivl_22508 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4037
  signal tmp_ivl_22510 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4037
  signal tmp_ivl_22515 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4037
  signal tmp_ivl_22517 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4037
  signal tmp_ivl_22519 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4037
  signal tmp_ivl_22521 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4037
  signal tmp_ivl_22526 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4038
  signal tmp_ivl_2253 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3017
  signal tmp_ivl_22531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4038
  signal tmp_ivl_22533 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4038
  signal tmp_ivl_22538 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4038
  signal tmp_ivl_22540 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4038
  signal tmp_ivl_22545 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4039
  signal tmp_ivl_2255 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3017
  signal tmp_ivl_22550 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4039
  signal tmp_ivl_22552 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4039
  signal tmp_ivl_22557 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4039
  signal tmp_ivl_22559 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4039
  signal tmp_ivl_22561 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4039
  signal tmp_ivl_22563 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4039
  signal tmp_ivl_22568 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4040
  signal tmp_ivl_2257 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3017
  signal tmp_ivl_22573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4040
  signal tmp_ivl_22575 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4040
  signal tmp_ivl_22580 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4040
  signal tmp_ivl_22582 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4040
  signal tmp_ivl_22588 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4041
  signal tmp_ivl_22589 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4041
  signal tmp_ivl_22594 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4041
  signal tmp_ivl_22597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4041
  signal tmp_ivl_22599 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4041
  signal tmp_ivl_22600 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4041
  signal tmp_ivl_22605 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4041
  signal tmp_ivl_22607 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4041
  signal tmp_ivl_22613 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4042
  signal tmp_ivl_22615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4042
  signal tmp_ivl_22616 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4042
  signal tmp_ivl_22621 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4042
  signal tmp_ivl_22623 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4042
  signal tmp_ivl_22628 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4042
  signal tmp_ivl_2263 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3018
  signal tmp_ivl_22630 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4042
  signal tmp_ivl_22635 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4043
  signal tmp_ivl_22640 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4043
  signal tmp_ivl_22642 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4043
  signal tmp_ivl_22647 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4043
  signal tmp_ivl_22649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4043
  signal tmp_ivl_2265 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3018
  signal tmp_ivl_22654 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4044
  signal tmp_ivl_22659 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4044
  signal tmp_ivl_2266 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3018
  signal tmp_ivl_22661 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4044
  signal tmp_ivl_22666 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4044
  signal tmp_ivl_22668 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4044
  signal tmp_ivl_22670 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4044
  signal tmp_ivl_22672 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4044
  signal tmp_ivl_22677 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4045
  signal tmp_ivl_22682 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4045
  signal tmp_ivl_22684 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4045
  signal tmp_ivl_22689 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4045
  signal tmp_ivl_22691 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4045
  signal tmp_ivl_22696 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4046
  signal tmp_ivl_227 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2947
  signal tmp_ivl_22701 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4046
  signal tmp_ivl_22703 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4046
  signal tmp_ivl_22708 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4046
  signal tmp_ivl_2271 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3018
  signal tmp_ivl_22710 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4046
  signal tmp_ivl_22712 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4046
  signal tmp_ivl_22714 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4046
  signal tmp_ivl_22719 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4047
  signal tmp_ivl_22724 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4047
  signal tmp_ivl_22726 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4047
  signal tmp_ivl_22731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4047
  signal tmp_ivl_22733 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4047
  signal tmp_ivl_22738 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4048
  signal tmp_ivl_2274 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3018
  signal tmp_ivl_22743 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4048
  signal tmp_ivl_22745 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4048
  signal tmp_ivl_22750 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4048
  signal tmp_ivl_22752 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4048
  signal tmp_ivl_22758 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4049
  signal tmp_ivl_2276 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3018
  signal tmp_ivl_22760 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4049
  signal tmp_ivl_22761 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4049
  signal tmp_ivl_22766 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4049
  signal tmp_ivl_22769 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4049
  signal tmp_ivl_2277 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3018
  signal tmp_ivl_22770 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4049
  signal tmp_ivl_22775 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4049
  signal tmp_ivl_22777 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4049
  signal tmp_ivl_22782 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4050
  signal tmp_ivl_22787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4050
  signal tmp_ivl_22789 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4050
  signal tmp_ivl_22794 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4050
  signal tmp_ivl_22796 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4050
  signal tmp_ivl_22801 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4051
  signal tmp_ivl_22806 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4051
  signal tmp_ivl_22808 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4051
  signal tmp_ivl_22813 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4051
  signal tmp_ivl_22815 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4051
  signal tmp_ivl_22817 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4051
  signal tmp_ivl_22819 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4051
  signal tmp_ivl_2282 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3018
  signal tmp_ivl_22824 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4052
  signal tmp_ivl_22829 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4052
  signal tmp_ivl_22831 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4052
  signal tmp_ivl_22836 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4052
  signal tmp_ivl_22838 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4052
  signal tmp_ivl_2284 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3018
  signal tmp_ivl_22843 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4053
  signal tmp_ivl_22848 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4053
  signal tmp_ivl_22850 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4053
  signal tmp_ivl_22855 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4053
  signal tmp_ivl_22857 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4053
  signal tmp_ivl_22859 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4053
  signal tmp_ivl_2286 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3018
  signal tmp_ivl_22861 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4053
  signal tmp_ivl_22866 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4054
  signal tmp_ivl_22871 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4054
  signal tmp_ivl_22873 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4054
  signal tmp_ivl_22878 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4054
  signal tmp_ivl_22880 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4054
  signal tmp_ivl_22886 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4055
  signal tmp_ivl_22888 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4055
  signal tmp_ivl_22889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4055
  signal tmp_ivl_22894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4055
  signal tmp_ivl_22896 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4055
  signal tmp_ivl_22901 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4055
  signal tmp_ivl_22903 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4055
  signal tmp_ivl_22908 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4056
  signal tmp_ivl_22913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4056
  signal tmp_ivl_22915 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4056
  signal tmp_ivl_2292 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3019
  signal tmp_ivl_22920 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4056
  signal tmp_ivl_22922 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4056
  signal tmp_ivl_22924 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4056
  signal tmp_ivl_22926 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4056
  signal tmp_ivl_22931 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4057
  signal tmp_ivl_22936 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4057
  signal tmp_ivl_22938 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4057
  signal tmp_ivl_2294 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3019
  signal tmp_ivl_22943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4057
  signal tmp_ivl_22945 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4057
  signal tmp_ivl_2295 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3019
  signal tmp_ivl_22950 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4058
  signal tmp_ivl_22955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4058
  signal tmp_ivl_22957 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4058
  signal tmp_ivl_22962 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4058
  signal tmp_ivl_22964 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4058
  signal tmp_ivl_22966 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4058
  signal tmp_ivl_22968 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4058
  signal tmp_ivl_22973 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4059
  signal tmp_ivl_22978 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4059
  signal tmp_ivl_22980 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4059
  signal tmp_ivl_22985 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4059
  signal tmp_ivl_22987 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4059
  signal tmp_ivl_22993 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4060
  signal tmp_ivl_22994 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4060
  signal tmp_ivl_22999 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4060
  signal tmp_ivl_2300 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3019
  signal tmp_ivl_23002 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4060
  signal tmp_ivl_23004 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4060
  signal tmp_ivl_23005 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4060
  signal tmp_ivl_23010 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4060
  signal tmp_ivl_23012 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4060
  signal tmp_ivl_23017 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4061
  signal tmp_ivl_23022 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4061
  signal tmp_ivl_23024 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4061
  signal tmp_ivl_23029 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4061
  signal tmp_ivl_2303 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3019
  signal tmp_ivl_23031 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4061
  signal tmp_ivl_23036 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4062
  signal tmp_ivl_23041 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4062
  signal tmp_ivl_23043 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4062
  signal tmp_ivl_23048 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4062
  signal tmp_ivl_2305 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3019
  signal tmp_ivl_23050 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4062
  signal tmp_ivl_23052 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4062
  signal tmp_ivl_23054 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4062
  signal tmp_ivl_23059 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4063
  signal tmp_ivl_2306 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3019
  signal tmp_ivl_23064 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4063
  signal tmp_ivl_23066 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4063
  signal tmp_ivl_23071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4063
  signal tmp_ivl_23073 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4063
  signal tmp_ivl_23078 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4064
  signal tmp_ivl_23083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4064
  signal tmp_ivl_23085 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4064
  signal tmp_ivl_23090 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4064
  signal tmp_ivl_23092 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4064
  signal tmp_ivl_23094 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4064
  signal tmp_ivl_23096 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4064
  signal tmp_ivl_23101 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4065
  signal tmp_ivl_23106 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4065
  signal tmp_ivl_23108 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4065
  signal tmp_ivl_2311 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3019
  signal tmp_ivl_23113 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4065
  signal tmp_ivl_23115 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4065
  signal tmp_ivl_23120 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4066
  signal tmp_ivl_23125 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4066
  signal tmp_ivl_23127 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4066
  signal tmp_ivl_2313 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3019
  signal tmp_ivl_23132 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4066
  signal tmp_ivl_23134 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4066
  signal tmp_ivl_23136 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4066
  signal tmp_ivl_23138 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4066
  signal tmp_ivl_23143 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4067
  signal tmp_ivl_23148 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4067
  signal tmp_ivl_2315 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3019
  signal tmp_ivl_23150 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4067
  signal tmp_ivl_23155 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4067
  signal tmp_ivl_23157 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4067
  signal tmp_ivl_23163 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4068
  signal tmp_ivl_23164 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4068
  signal tmp_ivl_23169 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4068
  signal tmp_ivl_23171 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4068
  signal tmp_ivl_23176 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4068
  signal tmp_ivl_23178 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4068
  signal tmp_ivl_23183 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4069
  signal tmp_ivl_23188 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4069
  signal tmp_ivl_23190 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4069
  signal tmp_ivl_23195 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4069
  signal tmp_ivl_23197 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4069
  signal tmp_ivl_23202 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4070
  signal tmp_ivl_23207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4070
  signal tmp_ivl_23209 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4070
  signal tmp_ivl_2321 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3020
  signal tmp_ivl_23214 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4070
  signal tmp_ivl_23216 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4070
  signal tmp_ivl_23218 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4070
  signal tmp_ivl_23220 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4070
  signal tmp_ivl_23225 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4071
  signal tmp_ivl_2323 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3020
  signal tmp_ivl_23230 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4071
  signal tmp_ivl_23232 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4071
  signal tmp_ivl_23237 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4071
  signal tmp_ivl_23239 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4071
  signal tmp_ivl_2324 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3020
  signal tmp_ivl_23244 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4072
  signal tmp_ivl_23249 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4072
  signal tmp_ivl_23251 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4072
  signal tmp_ivl_23256 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4072
  signal tmp_ivl_23258 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4072
  signal tmp_ivl_23260 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4072
  signal tmp_ivl_23262 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4072
  signal tmp_ivl_23267 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4073
  signal tmp_ivl_23272 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4073
  signal tmp_ivl_23274 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4073
  signal tmp_ivl_23279 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4073
  signal tmp_ivl_23281 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4073
  signal tmp_ivl_23287 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4074
  signal tmp_ivl_23288 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4074
  signal tmp_ivl_2329 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3020
  signal tmp_ivl_23293 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4074
  signal tmp_ivl_23296 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4074
  signal tmp_ivl_23298 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4074
  signal tmp_ivl_23299 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4074
  signal tmp_ivl_233 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2948
  signal tmp_ivl_23304 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4074
  signal tmp_ivl_23306 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4074
  signal tmp_ivl_23311 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4075
  signal tmp_ivl_23316 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4075
  signal tmp_ivl_23318 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4075
  signal tmp_ivl_2332 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3020
  signal tmp_ivl_23323 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4075
  signal tmp_ivl_23325 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4075
  signal tmp_ivl_23330 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4076
  signal tmp_ivl_23335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4076
  signal tmp_ivl_23337 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4076
  signal tmp_ivl_2334 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3020
  signal tmp_ivl_23342 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4076
  signal tmp_ivl_23344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4076
  signal tmp_ivl_23346 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4076
  signal tmp_ivl_23348 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4076
  signal tmp_ivl_2335 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3020
  signal tmp_ivl_23353 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4077
  signal tmp_ivl_23358 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4077
  signal tmp_ivl_23360 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4077
  signal tmp_ivl_23365 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4077
  signal tmp_ivl_23367 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4077
  signal tmp_ivl_23372 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4078
  signal tmp_ivl_23377 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4078
  signal tmp_ivl_23379 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4078
  signal tmp_ivl_23384 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4078
  signal tmp_ivl_23386 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4078
  signal tmp_ivl_23388 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4078
  signal tmp_ivl_23390 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4078
  signal tmp_ivl_23395 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4079
  signal tmp_ivl_2340 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3020
  signal tmp_ivl_23400 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4079
  signal tmp_ivl_23402 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4079
  signal tmp_ivl_23407 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4079
  signal tmp_ivl_23409 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4079
  signal tmp_ivl_23414 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4080
  signal tmp_ivl_23419 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4080
  signal tmp_ivl_2342 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3020
  signal tmp_ivl_23421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4080
  signal tmp_ivl_23426 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4080
  signal tmp_ivl_23428 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4080
  signal tmp_ivl_23430 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4080
  signal tmp_ivl_23432 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4080
  signal tmp_ivl_23437 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4081
  signal tmp_ivl_2344 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3020
  signal tmp_ivl_23442 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4081
  signal tmp_ivl_23444 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4081
  signal tmp_ivl_23449 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4081
  signal tmp_ivl_23451 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4081
  signal tmp_ivl_23457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4082
  signal tmp_ivl_23458 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4082
  signal tmp_ivl_23463 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4082
  signal tmp_ivl_23466 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4082
  signal tmp_ivl_23468 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4082
  signal tmp_ivl_23469 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4082
  signal tmp_ivl_23474 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4082
  signal tmp_ivl_23476 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4082
  signal tmp_ivl_23482 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4083
  signal tmp_ivl_23484 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4083
  signal tmp_ivl_23485 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4083
  signal tmp_ivl_23490 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4083
  signal tmp_ivl_23492 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4083
  signal tmp_ivl_23497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4083
  signal tmp_ivl_23499 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4083
  signal tmp_ivl_235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2948
  signal tmp_ivl_2350 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3021
  signal tmp_ivl_23504 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4084
  signal tmp_ivl_23509 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4084
  signal tmp_ivl_23511 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4084
  signal tmp_ivl_23516 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4084
  signal tmp_ivl_23518 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4084
  signal tmp_ivl_2352 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3021
  signal tmp_ivl_23523 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4085
  signal tmp_ivl_23528 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4085
  signal tmp_ivl_2353 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3021
  signal tmp_ivl_23530 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4085
  signal tmp_ivl_23535 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4085
  signal tmp_ivl_23537 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4085
  signal tmp_ivl_23539 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4085
  signal tmp_ivl_23541 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4085
  signal tmp_ivl_23546 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4086
  signal tmp_ivl_23551 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4086
  signal tmp_ivl_23553 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4086
  signal tmp_ivl_23558 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4086
  signal tmp_ivl_23560 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4086
  signal tmp_ivl_23565 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4087
  signal tmp_ivl_23570 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4087
  signal tmp_ivl_23572 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4087
  signal tmp_ivl_23577 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4087
  signal tmp_ivl_23579 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4087
  signal tmp_ivl_2358 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3021
  signal tmp_ivl_23581 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4087
  signal tmp_ivl_23583 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4087
  signal tmp_ivl_23588 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4088
  signal tmp_ivl_23593 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4088
  signal tmp_ivl_23595 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4088
  signal tmp_ivl_236 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2948
  signal tmp_ivl_23600 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4088
  signal tmp_ivl_23602 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4088
  signal tmp_ivl_23607 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4089
  signal tmp_ivl_2361 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3021
  signal tmp_ivl_23612 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4089
  signal tmp_ivl_23614 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4089
  signal tmp_ivl_23619 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4089
  signal tmp_ivl_23621 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4089
  signal tmp_ivl_23623 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4089
  signal tmp_ivl_23625 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4089
  signal tmp_ivl_2363 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3021
  signal tmp_ivl_23630 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4090
  signal tmp_ivl_23635 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4090
  signal tmp_ivl_23637 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4090
  signal tmp_ivl_2364 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3021
  signal tmp_ivl_23642 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4090
  signal tmp_ivl_23644 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4090
  signal tmp_ivl_23650 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4091
  signal tmp_ivl_23652 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4091
  signal tmp_ivl_23653 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4091
  signal tmp_ivl_23658 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4091
  signal tmp_ivl_23661 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4091
  signal tmp_ivl_23662 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4091
  signal tmp_ivl_23667 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4091
  signal tmp_ivl_23669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4091
  signal tmp_ivl_23674 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4092
  signal tmp_ivl_23679 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4092
  signal tmp_ivl_23681 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4092
  signal tmp_ivl_23686 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4092
  signal tmp_ivl_23688 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4092
  signal tmp_ivl_2369 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3021
  signal tmp_ivl_23693 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4093
  signal tmp_ivl_23698 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4093
  signal tmp_ivl_23700 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4093
  signal tmp_ivl_23705 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4093
  signal tmp_ivl_23707 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4093
  signal tmp_ivl_23709 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4093
  signal tmp_ivl_2371 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3021
  signal tmp_ivl_23711 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4093
  signal tmp_ivl_23716 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4094
  signal tmp_ivl_23721 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4094
  signal tmp_ivl_23723 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4094
  signal tmp_ivl_23728 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4094
  signal tmp_ivl_2373 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3021
  signal tmp_ivl_23730 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4094
  signal tmp_ivl_23735 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4095
  signal tmp_ivl_23740 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4095
  signal tmp_ivl_23742 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4095
  signal tmp_ivl_23747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4095
  signal tmp_ivl_23749 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4095
  signal tmp_ivl_23751 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4095
  signal tmp_ivl_23753 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4095
  signal tmp_ivl_23758 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4096
  signal tmp_ivl_23763 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4096
  signal tmp_ivl_23765 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4096
  signal tmp_ivl_23770 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4096
  signal tmp_ivl_23772 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4096
  signal tmp_ivl_23777 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4097
  signal tmp_ivl_23782 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4097
  signal tmp_ivl_23784 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4097
  signal tmp_ivl_23789 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4097
  signal tmp_ivl_2379 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3022
  signal tmp_ivl_23791 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4097
  signal tmp_ivl_23793 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4097
  signal tmp_ivl_23795 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4097
  signal tmp_ivl_23800 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4098
  signal tmp_ivl_23805 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4098
  signal tmp_ivl_23807 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4098
  signal tmp_ivl_2381 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3022
  signal tmp_ivl_23812 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4098
  signal tmp_ivl_23814 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4098
  signal tmp_ivl_2382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3022
  signal tmp_ivl_23820 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4099
  signal tmp_ivl_23822 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4099
  signal tmp_ivl_23823 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4099
  signal tmp_ivl_23828 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4099
  signal tmp_ivl_23830 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4099
  signal tmp_ivl_23835 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4099
  signal tmp_ivl_23837 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4099
  signal tmp_ivl_23842 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4100
  signal tmp_ivl_23847 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4100
  signal tmp_ivl_23849 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4100
  signal tmp_ivl_23854 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4100
  signal tmp_ivl_23856 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4100
  signal tmp_ivl_23858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4100
  signal tmp_ivl_23860 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4100
  signal tmp_ivl_23865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4101
  signal tmp_ivl_2387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3022
  signal tmp_ivl_23870 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4101
  signal tmp_ivl_23872 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4101
  signal tmp_ivl_23877 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4101
  signal tmp_ivl_23879 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4101
  signal tmp_ivl_23884 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4102
  signal tmp_ivl_23889 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4102
  signal tmp_ivl_23891 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4102
  signal tmp_ivl_23896 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4102
  signal tmp_ivl_23898 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4102
  signal tmp_ivl_2390 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3022
  signal tmp_ivl_23900 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4102
  signal tmp_ivl_23902 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4102
  signal tmp_ivl_23907 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4103
  signal tmp_ivl_23912 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4103
  signal tmp_ivl_23914 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4103
  signal tmp_ivl_23919 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4103
  signal tmp_ivl_2392 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3022
  signal tmp_ivl_23921 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4103
  signal tmp_ivl_23926 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4104
  signal tmp_ivl_2393 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3022
  signal tmp_ivl_23931 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4104
  signal tmp_ivl_23933 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4104
  signal tmp_ivl_23938 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4104
  signal tmp_ivl_23940 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4104
  signal tmp_ivl_23942 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4104
  signal tmp_ivl_23944 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4104
  signal tmp_ivl_23949 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4105
  signal tmp_ivl_23954 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4105
  signal tmp_ivl_23956 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4105
  signal tmp_ivl_23961 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4105
  signal tmp_ivl_23963 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4105
  signal tmp_ivl_23969 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4106
  signal tmp_ivl_23970 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4106
  signal tmp_ivl_23975 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4106
  signal tmp_ivl_23978 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4106
  signal tmp_ivl_2398 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3022
  signal tmp_ivl_23980 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4106
  signal tmp_ivl_23981 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4106
  signal tmp_ivl_23986 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4106
  signal tmp_ivl_23988 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4106
  signal tmp_ivl_23993 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4107
  signal tmp_ivl_23998 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4107
  signal tmp_ivl_24 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2940
  signal tmp_ivl_2400 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3022
  signal tmp_ivl_24000 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4107
  signal tmp_ivl_24005 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4107
  signal tmp_ivl_24007 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4107
  signal tmp_ivl_24012 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4108
  signal tmp_ivl_24017 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4108
  signal tmp_ivl_24019 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4108
  signal tmp_ivl_2402 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3022
  signal tmp_ivl_24024 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4108
  signal tmp_ivl_24026 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4108
  signal tmp_ivl_24028 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4108
  signal tmp_ivl_24030 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4108
  signal tmp_ivl_24035 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4109
  signal tmp_ivl_24040 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4109
  signal tmp_ivl_24042 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4109
  signal tmp_ivl_24047 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4109
  signal tmp_ivl_24049 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4109
  signal tmp_ivl_24054 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4110
  signal tmp_ivl_24059 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4110
  signal tmp_ivl_24061 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4110
  signal tmp_ivl_24066 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4110
  signal tmp_ivl_24068 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4110
  signal tmp_ivl_24070 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4110
  signal tmp_ivl_24072 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4110
  signal tmp_ivl_24077 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4111
  signal tmp_ivl_2408 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3023
  signal tmp_ivl_24082 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4111
  signal tmp_ivl_24084 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4111
  signal tmp_ivl_24089 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4111
  signal tmp_ivl_24091 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4111
  signal tmp_ivl_24097 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4112
  signal tmp_ivl_24098 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4112
  signal tmp_ivl_241 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2948
  signal tmp_ivl_2410 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3023
  signal tmp_ivl_24103 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4112
  signal tmp_ivl_24106 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4112
  signal tmp_ivl_24108 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4112
  signal tmp_ivl_24109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4112
  signal tmp_ivl_2411 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3023
  signal tmp_ivl_24114 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4112
  signal tmp_ivl_24116 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4112
  signal tmp_ivl_24122 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4113
  signal tmp_ivl_24124 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4113
  signal tmp_ivl_24125 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4113
  signal tmp_ivl_24130 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4113
  signal tmp_ivl_24132 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4113
  signal tmp_ivl_24137 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4113
  signal tmp_ivl_24139 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4113
  signal tmp_ivl_24144 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4114
  signal tmp_ivl_24149 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4114
  signal tmp_ivl_24151 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4114
  signal tmp_ivl_24156 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4114
  signal tmp_ivl_24158 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4114
  signal tmp_ivl_2416 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3023
  signal tmp_ivl_24163 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4115
  signal tmp_ivl_24168 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4115
  signal tmp_ivl_24170 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4115
  signal tmp_ivl_24175 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4115
  signal tmp_ivl_24177 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4115
  signal tmp_ivl_24179 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4115
  signal tmp_ivl_24181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4115
  signal tmp_ivl_24186 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4116
  signal tmp_ivl_2419 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3023
  signal tmp_ivl_24191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4116
  signal tmp_ivl_24193 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4116
  signal tmp_ivl_24198 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4116
  signal tmp_ivl_24200 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4116
  signal tmp_ivl_24205 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4117
  signal tmp_ivl_2421 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3023
  signal tmp_ivl_24210 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4117
  signal tmp_ivl_24212 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4117
  signal tmp_ivl_24217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4117
  signal tmp_ivl_24219 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4117
  signal tmp_ivl_2422 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3023
  signal tmp_ivl_24221 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4117
  signal tmp_ivl_24223 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4117
  signal tmp_ivl_24228 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4118
  signal tmp_ivl_24233 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4118
  signal tmp_ivl_24235 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4118
  signal tmp_ivl_24240 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4118
  signal tmp_ivl_24242 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4118
  signal tmp_ivl_24248 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4119
  signal tmp_ivl_24250 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4119
  signal tmp_ivl_24251 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4119
  signal tmp_ivl_24256 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4119
  signal tmp_ivl_24259 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4119
  signal tmp_ivl_24260 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4119
  signal tmp_ivl_24265 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4119
  signal tmp_ivl_24267 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4119
  signal tmp_ivl_2427 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3023
  signal tmp_ivl_24272 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4120
  signal tmp_ivl_24277 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4120
  signal tmp_ivl_24279 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4120
  signal tmp_ivl_24284 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4120
  signal tmp_ivl_24286 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4120
  signal tmp_ivl_2429 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3023
  signal tmp_ivl_24291 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4121
  signal tmp_ivl_24296 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4121
  signal tmp_ivl_24298 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4121
  signal tmp_ivl_24303 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4121
  signal tmp_ivl_24305 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4121
  signal tmp_ivl_24307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4121
  signal tmp_ivl_24309 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4121
  signal tmp_ivl_2431 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3023
  signal tmp_ivl_24314 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4122
  signal tmp_ivl_24319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4122
  signal tmp_ivl_24321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4122
  signal tmp_ivl_24326 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4122
  signal tmp_ivl_24328 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4122
  signal tmp_ivl_24333 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4123
  signal tmp_ivl_24338 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4123
  signal tmp_ivl_24340 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4123
  signal tmp_ivl_24345 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4123
  signal tmp_ivl_24347 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4123
  signal tmp_ivl_24349 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4123
  signal tmp_ivl_24351 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4123
  signal tmp_ivl_24356 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4124
  signal tmp_ivl_24361 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4124
  signal tmp_ivl_24363 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4124
  signal tmp_ivl_24368 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4124
  signal tmp_ivl_2437 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3024
  signal tmp_ivl_24370 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4124
  signal tmp_ivl_24375 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4125
  signal tmp_ivl_24380 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4125
  signal tmp_ivl_24382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4125
  signal tmp_ivl_24387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4125
  signal tmp_ivl_24389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4125
  signal tmp_ivl_2439 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3024
  signal tmp_ivl_24391 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4125
  signal tmp_ivl_24393 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4125
  signal tmp_ivl_24398 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4126
  signal tmp_ivl_244 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2948
  signal tmp_ivl_2440 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3024
  signal tmp_ivl_24403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4126
  signal tmp_ivl_24405 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4126
  signal tmp_ivl_24410 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4126
  signal tmp_ivl_24412 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4126
  signal tmp_ivl_24418 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4127
  signal tmp_ivl_24420 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4127
  signal tmp_ivl_24421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4127
  signal tmp_ivl_24426 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4127
  signal tmp_ivl_24428 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4127
  signal tmp_ivl_24433 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4127
  signal tmp_ivl_24435 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4127
  signal tmp_ivl_24440 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4128
  signal tmp_ivl_24445 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4128
  signal tmp_ivl_24447 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4128
  signal tmp_ivl_2445 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3024
  signal tmp_ivl_24452 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4128
  signal tmp_ivl_24454 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4128
  signal tmp_ivl_24456 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4128
  signal tmp_ivl_24458 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4128
  signal tmp_ivl_24463 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4129
  signal tmp_ivl_24468 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4129
  signal tmp_ivl_24470 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4129
  signal tmp_ivl_24475 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4129
  signal tmp_ivl_24477 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4129
  signal tmp_ivl_2448 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3024
  signal tmp_ivl_24482 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4130
  signal tmp_ivl_24487 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4130
  signal tmp_ivl_24489 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4130
  signal tmp_ivl_24494 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4130
  signal tmp_ivl_24496 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4130
  signal tmp_ivl_24498 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4130
  signal tmp_ivl_2450 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3024
  signal tmp_ivl_24500 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4130
  signal tmp_ivl_24505 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4131
  signal tmp_ivl_2451 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3024
  signal tmp_ivl_24510 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4131
  signal tmp_ivl_24512 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4131
  signal tmp_ivl_24517 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4131
  signal tmp_ivl_24519 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4131
  signal tmp_ivl_24525 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4132
  signal tmp_ivl_24526 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4132
  signal tmp_ivl_24531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4132
  signal tmp_ivl_24534 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4132
  signal tmp_ivl_24536 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4132
  signal tmp_ivl_24537 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4132
  signal tmp_ivl_24542 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4132
  signal tmp_ivl_24544 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4132
  signal tmp_ivl_24549 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4133
  signal tmp_ivl_24554 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4133
  signal tmp_ivl_24556 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4133
  signal tmp_ivl_2456 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3024
  signal tmp_ivl_24561 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4133
  signal tmp_ivl_24563 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4133
  signal tmp_ivl_24568 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4134
  signal tmp_ivl_24573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4134
  signal tmp_ivl_24575 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4134
  signal tmp_ivl_2458 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3024
  signal tmp_ivl_24580 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4134
  signal tmp_ivl_24582 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4134
  signal tmp_ivl_24584 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4134
  signal tmp_ivl_24586 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4134
  signal tmp_ivl_24591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4135
  signal tmp_ivl_24596 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4135
  signal tmp_ivl_24598 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4135
  signal tmp_ivl_246 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2948
  signal tmp_ivl_2460 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3024
  signal tmp_ivl_24603 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4135
  signal tmp_ivl_24605 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4135
  signal tmp_ivl_24610 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4136
  signal tmp_ivl_24615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4136
  signal tmp_ivl_24617 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4136
  signal tmp_ivl_24622 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4136
  signal tmp_ivl_24624 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4136
  signal tmp_ivl_24626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4136
  signal tmp_ivl_24628 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4136
  signal tmp_ivl_24633 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4137
  signal tmp_ivl_24638 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4137
  signal tmp_ivl_24640 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4137
  signal tmp_ivl_24645 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4137
  signal tmp_ivl_24647 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4137
  signal tmp_ivl_24653 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4138
  signal tmp_ivl_24654 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4138
  signal tmp_ivl_24659 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4138
  signal tmp_ivl_2466 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3025
  signal tmp_ivl_24662 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4138
  signal tmp_ivl_24664 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4138
  signal tmp_ivl_24665 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4138
  signal tmp_ivl_24670 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4138
  signal tmp_ivl_24672 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4138
  signal tmp_ivl_24678 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4139
  signal tmp_ivl_2468 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3025
  signal tmp_ivl_24680 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4139
  signal tmp_ivl_24681 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4139
  signal tmp_ivl_24686 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4139
  signal tmp_ivl_24688 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4139
  signal tmp_ivl_2469 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3025
  signal tmp_ivl_24693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4139
  signal tmp_ivl_24695 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4139
  signal tmp_ivl_247 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2948
  signal tmp_ivl_24700 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4140
  signal tmp_ivl_24705 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4140
  signal tmp_ivl_24707 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4140
  signal tmp_ivl_24712 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4140
  signal tmp_ivl_24714 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4140
  signal tmp_ivl_24719 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4141
  signal tmp_ivl_24724 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4141
  signal tmp_ivl_24726 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4141
  signal tmp_ivl_24731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4141
  signal tmp_ivl_24733 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4141
  signal tmp_ivl_24735 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4141
  signal tmp_ivl_24737 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4141
  signal tmp_ivl_2474 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3025
  signal tmp_ivl_24742 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4142
  signal tmp_ivl_24747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4142
  signal tmp_ivl_24749 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4142
  signal tmp_ivl_24754 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4142
  signal tmp_ivl_24756 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4142
  signal tmp_ivl_24761 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4143
  signal tmp_ivl_24766 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4143
  signal tmp_ivl_24768 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4143
  signal tmp_ivl_2477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3025
  signal tmp_ivl_24773 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4143
  signal tmp_ivl_24775 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4143
  signal tmp_ivl_24777 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4143
  signal tmp_ivl_24779 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4143
  signal tmp_ivl_24784 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4144
  signal tmp_ivl_24789 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4144
  signal tmp_ivl_2479 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3025
  signal tmp_ivl_24791 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4144
  signal tmp_ivl_24796 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4144
  signal tmp_ivl_24798 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4144
  signal tmp_ivl_2480 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3025
  signal tmp_ivl_24804 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4145
  signal tmp_ivl_24805 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4145
  signal tmp_ivl_24810 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4145
  signal tmp_ivl_24813 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4145
  signal tmp_ivl_24815 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4145
  signal tmp_ivl_24816 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4145
  signal tmp_ivl_24821 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4145
  signal tmp_ivl_24823 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4145
  signal tmp_ivl_24828 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4146
  signal tmp_ivl_24833 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4146
  signal tmp_ivl_24835 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4146
  signal tmp_ivl_24840 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4146
  signal tmp_ivl_24842 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4146
  signal tmp_ivl_24847 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4147
  signal tmp_ivl_2485 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3025
  signal tmp_ivl_24852 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4147
  signal tmp_ivl_24854 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4147
  signal tmp_ivl_24859 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4147
  signal tmp_ivl_24861 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4147
  signal tmp_ivl_24863 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4147
  signal tmp_ivl_24865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4147
  signal tmp_ivl_2487 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3025
  signal tmp_ivl_24870 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4148
  signal tmp_ivl_24875 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4148
  signal tmp_ivl_24877 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4148
  signal tmp_ivl_24882 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4148
  signal tmp_ivl_24884 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4148
  signal tmp_ivl_24889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4149
  signal tmp_ivl_2489 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3025
  signal tmp_ivl_24894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4149
  signal tmp_ivl_24896 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4149
  signal tmp_ivl_24901 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4149
  signal tmp_ivl_24903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4149
  signal tmp_ivl_24905 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4149
  signal tmp_ivl_24907 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4149
  signal tmp_ivl_24912 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4150
  signal tmp_ivl_24917 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4150
  signal tmp_ivl_24919 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4150
  signal tmp_ivl_24924 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4150
  signal tmp_ivl_24926 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4150
  signal tmp_ivl_24931 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4151
  signal tmp_ivl_24936 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4151
  signal tmp_ivl_24938 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4151
  signal tmp_ivl_24943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4151
  signal tmp_ivl_24945 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4151
  signal tmp_ivl_24947 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4151
  signal tmp_ivl_24949 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4151
  signal tmp_ivl_2495 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3026
  signal tmp_ivl_24954 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4152
  signal tmp_ivl_24959 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4152
  signal tmp_ivl_24961 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4152
  signal tmp_ivl_24966 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4152
  signal tmp_ivl_24968 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4152
  signal tmp_ivl_2497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3026
  signal tmp_ivl_24974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4153
  signal tmp_ivl_24975 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4153
  signal tmp_ivl_2498 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3026
  signal tmp_ivl_24980 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4153
  signal tmp_ivl_24983 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4153
  signal tmp_ivl_24985 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4153
  signal tmp_ivl_24986 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4153
  signal tmp_ivl_24991 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4153
  signal tmp_ivl_24993 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4153
  signal tmp_ivl_24999 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4154
  signal tmp_ivl_25001 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4154
  signal tmp_ivl_25002 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4154
  signal tmp_ivl_25007 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4154
  signal tmp_ivl_25009 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4154
  signal tmp_ivl_25014 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4154
  signal tmp_ivl_25016 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4154
  signal tmp_ivl_25021 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4155
  signal tmp_ivl_25026 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4155
  signal tmp_ivl_25028 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4155
  signal tmp_ivl_2503 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3026
  signal tmp_ivl_25033 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4155
  signal tmp_ivl_25035 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4155
  signal tmp_ivl_25040 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4156
  signal tmp_ivl_25045 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4156
  signal tmp_ivl_25047 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4156
  signal tmp_ivl_25052 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4156
  signal tmp_ivl_25054 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4156
  signal tmp_ivl_25056 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4156
  signal tmp_ivl_25058 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4156
  signal tmp_ivl_2506 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3026
  signal tmp_ivl_25063 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4157
  signal tmp_ivl_25068 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4157
  signal tmp_ivl_25070 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4157
  signal tmp_ivl_25075 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4157
  signal tmp_ivl_25077 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4157
  signal tmp_ivl_2508 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3026
  signal tmp_ivl_25082 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4158
  signal tmp_ivl_25087 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4158
  signal tmp_ivl_25089 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4158
  signal tmp_ivl_2509 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3026
  signal tmp_ivl_25094 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4158
  signal tmp_ivl_25096 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4158
  signal tmp_ivl_25098 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4158
  signal tmp_ivl_25100 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4158
  signal tmp_ivl_25105 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4159
  signal tmp_ivl_25110 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4159
  signal tmp_ivl_25112 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4159
  signal tmp_ivl_25117 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4159
  signal tmp_ivl_25119 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4159
  signal tmp_ivl_25124 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4160
  signal tmp_ivl_25129 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4160
  signal tmp_ivl_25131 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4160
  signal tmp_ivl_25136 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4160
  signal tmp_ivl_25138 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4160
  signal tmp_ivl_2514 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3026
  signal tmp_ivl_25140 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4160
  signal tmp_ivl_25142 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4160
  signal tmp_ivl_25147 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4161
  signal tmp_ivl_25152 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4161
  signal tmp_ivl_25154 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4161
  signal tmp_ivl_25159 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4161
  signal tmp_ivl_2516 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3026
  signal tmp_ivl_25161 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4161
  signal tmp_ivl_25167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4162
  signal tmp_ivl_25169 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4162
  signal tmp_ivl_25170 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4162
  signal tmp_ivl_25175 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4162
  signal tmp_ivl_25178 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4162
  signal tmp_ivl_25179 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4162
  signal tmp_ivl_2518 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3026
  signal tmp_ivl_25184 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4162
  signal tmp_ivl_25186 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4162
  signal tmp_ivl_25191 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4163
  signal tmp_ivl_25196 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4163
  signal tmp_ivl_25198 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4163
  signal tmp_ivl_252 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2948
  signal tmp_ivl_25203 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4163
  signal tmp_ivl_25205 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4163
  signal tmp_ivl_25210 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4164
  signal tmp_ivl_25215 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4164
  signal tmp_ivl_25217 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4164
  signal tmp_ivl_25222 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4164
  signal tmp_ivl_25224 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4164
  signal tmp_ivl_25226 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4164
  signal tmp_ivl_25228 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4164
  signal tmp_ivl_25233 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4165
  signal tmp_ivl_25238 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4165
  signal tmp_ivl_2524 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3027
  signal tmp_ivl_25240 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4165
  signal tmp_ivl_25245 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4165
  signal tmp_ivl_25247 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4165
  signal tmp_ivl_25252 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4166
  signal tmp_ivl_25257 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4166
  signal tmp_ivl_25259 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4166
  signal tmp_ivl_2526 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3027
  signal tmp_ivl_25264 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4166
  signal tmp_ivl_25266 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4166
  signal tmp_ivl_25268 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4166
  signal tmp_ivl_2527 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3027
  signal tmp_ivl_25270 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4166
  signal tmp_ivl_25275 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4167
  signal tmp_ivl_25280 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4167
  signal tmp_ivl_25282 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4167
  signal tmp_ivl_25287 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4167
  signal tmp_ivl_25289 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4167
  signal tmp_ivl_25294 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4168
  signal tmp_ivl_25299 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4168
  signal tmp_ivl_25301 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4168
  signal tmp_ivl_25306 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4168
  signal tmp_ivl_25308 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4168
  signal tmp_ivl_25310 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4168
  signal tmp_ivl_25312 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4168
  signal tmp_ivl_25317 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4169
  signal tmp_ivl_2532 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3027
  signal tmp_ivl_25322 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4169
  signal tmp_ivl_25324 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4169
  signal tmp_ivl_25329 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4169
  signal tmp_ivl_25331 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4169
  signal tmp_ivl_25337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4170
  signal tmp_ivl_25339 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4170
  signal tmp_ivl_25340 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4170
  signal tmp_ivl_25345 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4170
  signal tmp_ivl_25347 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4170
  signal tmp_ivl_2535 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3027
  signal tmp_ivl_25352 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4170
  signal tmp_ivl_25354 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4170
  signal tmp_ivl_25359 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4171
  signal tmp_ivl_25364 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4171
  signal tmp_ivl_25366 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4171
  signal tmp_ivl_2537 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3027
  signal tmp_ivl_25371 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4171
  signal tmp_ivl_25373 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4171
  signal tmp_ivl_25375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4171
  signal tmp_ivl_25377 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4171
  signal tmp_ivl_2538 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3027
  signal tmp_ivl_25382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4172
  signal tmp_ivl_25387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4172
  signal tmp_ivl_25389 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4172
  signal tmp_ivl_25394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4172
  signal tmp_ivl_25396 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4172
  signal tmp_ivl_254 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2948
  signal tmp_ivl_25401 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4173
  signal tmp_ivl_25406 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4173
  signal tmp_ivl_25408 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4173
  signal tmp_ivl_25413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4173
  signal tmp_ivl_25415 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4173
  signal tmp_ivl_25417 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4173
  signal tmp_ivl_25419 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4173
  signal tmp_ivl_25424 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4174
  signal tmp_ivl_25429 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4174
  signal tmp_ivl_2543 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3027
  signal tmp_ivl_25431 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4174
  signal tmp_ivl_25436 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4174
  signal tmp_ivl_25438 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4174
  signal tmp_ivl_25443 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4175
  signal tmp_ivl_25448 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4175
  signal tmp_ivl_2545 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3027
  signal tmp_ivl_25450 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4175
  signal tmp_ivl_25455 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4175
  signal tmp_ivl_25457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4175
  signal tmp_ivl_25459 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4175
  signal tmp_ivl_25461 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4175
  signal tmp_ivl_25466 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4176
  signal tmp_ivl_2547 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3027
  signal tmp_ivl_25471 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4176
  signal tmp_ivl_25474 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4176
  signal tmp_ivl_25475 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4176
  signal tmp_ivl_25480 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4176
  signal tmp_ivl_25482 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4176
  signal tmp_ivl_25488 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4177
  signal tmp_ivl_25489 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4177
  signal tmp_ivl_25494 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4177
  signal tmp_ivl_25497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4177
  signal tmp_ivl_25499 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4177
  signal tmp_ivl_25500 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4177
  signal tmp_ivl_25505 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4177
  signal tmp_ivl_25507 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4177
  signal tmp_ivl_25512 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4178
  signal tmp_ivl_25517 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4178
  signal tmp_ivl_25519 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4178
  signal tmp_ivl_25524 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4178
  signal tmp_ivl_25526 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4178
  signal tmp_ivl_2553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3028
  signal tmp_ivl_25531 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4179
  signal tmp_ivl_25536 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4179
  signal tmp_ivl_25539 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4179
  signal tmp_ivl_25540 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4179
  signal tmp_ivl_25545 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4179
  signal tmp_ivl_25547 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4179
  signal tmp_ivl_2555 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3028
  signal tmp_ivl_25553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4180
  signal tmp_ivl_25554 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4180
  signal tmp_ivl_25559 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4180
  signal tmp_ivl_2556 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3028
  signal tmp_ivl_25562 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4180
  signal tmp_ivl_25564 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4180
  signal tmp_ivl_25565 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4180
  signal tmp_ivl_25570 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4180
  signal tmp_ivl_25572 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4180
  signal tmp_ivl_25577 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4181
  signal tmp_ivl_25582 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4181
  signal tmp_ivl_25584 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4181
  signal tmp_ivl_25589 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4181
  signal tmp_ivl_25591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4181
  signal tmp_ivl_25596 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4182
  signal tmp_ivl_256 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2948
  signal tmp_ivl_25601 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4182
  signal tmp_ivl_25603 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4182
  signal tmp_ivl_25608 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4182
  signal tmp_ivl_2561 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3028
  signal tmp_ivl_25610 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4182
  signal tmp_ivl_25615 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4183
  signal tmp_ivl_25620 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4183
  signal tmp_ivl_25623 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4183
  signal tmp_ivl_25624 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4183
  signal tmp_ivl_25629 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4183
  signal tmp_ivl_25631 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4183
  signal tmp_ivl_25637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4184
  signal tmp_ivl_25638 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4184
  signal tmp_ivl_2564 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3028
  signal tmp_ivl_25643 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4184
  signal tmp_ivl_25646 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4184
  signal tmp_ivl_25648 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4184
  signal tmp_ivl_25649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4184
  signal tmp_ivl_25654 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4184
  signal tmp_ivl_25656 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4184
  signal tmp_ivl_2566 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3028
  signal tmp_ivl_25661 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4185
  signal tmp_ivl_25666 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4185
  signal tmp_ivl_25668 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4185
  signal tmp_ivl_2567 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3028
  signal tmp_ivl_25673 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4185
  signal tmp_ivl_25675 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4185
  signal tmp_ivl_25680 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4186
  signal tmp_ivl_25685 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4186
  signal tmp_ivl_25687 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4186
  signal tmp_ivl_25692 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4186
  signal tmp_ivl_25694 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4186
  signal tmp_ivl_25696 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4186
  signal tmp_ivl_25698 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4186
  signal tmp_ivl_25703 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4187
  signal tmp_ivl_25708 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4187
  signal tmp_ivl_25711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4187
  signal tmp_ivl_25712 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4187
  signal tmp_ivl_25717 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4187
  signal tmp_ivl_25719 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4187
  signal tmp_ivl_2572 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3028
  signal tmp_ivl_25725 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4188
  signal tmp_ivl_25726 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4188
  signal tmp_ivl_25731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4188
  signal tmp_ivl_25734 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4188
  signal tmp_ivl_25736 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4188
  signal tmp_ivl_25737 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4188
  signal tmp_ivl_2574 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3028
  signal tmp_ivl_25742 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4188
  signal tmp_ivl_25744 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4188
  signal tmp_ivl_25749 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4189
  signal tmp_ivl_25754 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4189
  signal tmp_ivl_25756 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4189
  signal tmp_ivl_2576 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3028
  signal tmp_ivl_25761 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4189
  signal tmp_ivl_25763 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4189
  signal tmp_ivl_25768 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4190
  signal tmp_ivl_25773 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4190
  signal tmp_ivl_25776 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4190
  signal tmp_ivl_25777 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4190
  signal tmp_ivl_25782 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4190
  signal tmp_ivl_25784 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4190
  signal tmp_ivl_25790 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4191
  signal tmp_ivl_25791 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4191
  signal tmp_ivl_25796 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4191
  signal tmp_ivl_25799 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4191
  signal tmp_ivl_25801 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4191
  signal tmp_ivl_25802 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4191
  signal tmp_ivl_25807 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4191
  signal tmp_ivl_25809 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4191
  signal tmp_ivl_25814 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4192
  signal tmp_ivl_25819 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4192
  signal tmp_ivl_2582 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3029
  signal tmp_ivl_25821 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4192
  signal tmp_ivl_25826 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4192
  signal tmp_ivl_25828 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4192
  signal tmp_ivl_25833 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4193
  signal tmp_ivl_25838 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4193
  signal tmp_ivl_2584 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3029
  signal tmp_ivl_25840 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4193
  signal tmp_ivl_25845 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4193
  signal tmp_ivl_25847 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4193
  signal tmp_ivl_2585 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3029
  signal tmp_ivl_25852 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4194
  signal tmp_ivl_25857 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4194
  signal tmp_ivl_25860 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4194
  signal tmp_ivl_25861 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4194
  signal tmp_ivl_25866 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4194
  signal tmp_ivl_25868 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4194
  signal tmp_ivl_25874 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4195
  signal tmp_ivl_25875 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4195
  signal tmp_ivl_25880 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4195
  signal tmp_ivl_25883 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4195
  signal tmp_ivl_25885 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4195
  signal tmp_ivl_25886 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4195
  signal tmp_ivl_25891 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4195
  signal tmp_ivl_25893 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4195
  signal tmp_ivl_25898 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4196
  signal tmp_ivl_2590 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3029
  signal tmp_ivl_25903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4196
  signal tmp_ivl_25905 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4196
  signal tmp_ivl_25910 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4196
  signal tmp_ivl_25912 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4196
  signal tmp_ivl_25917 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4197
  signal tmp_ivl_25922 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4197
  signal tmp_ivl_25924 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4197
  signal tmp_ivl_25929 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4197
  signal tmp_ivl_2593 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3029
  signal tmp_ivl_25931 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4197
  signal tmp_ivl_25933 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4197
  signal tmp_ivl_25935 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4197
  signal tmp_ivl_25940 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4198
  signal tmp_ivl_25945 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4198
  signal tmp_ivl_25948 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4198
  signal tmp_ivl_25949 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4198
  signal tmp_ivl_2595 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3029
  signal tmp_ivl_25954 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4198
  signal tmp_ivl_25956 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4198
  signal tmp_ivl_2596 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3029
  signal tmp_ivl_25962 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4199
  signal tmp_ivl_25963 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4199
  signal tmp_ivl_25968 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4199
  signal tmp_ivl_25971 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4199
  signal tmp_ivl_25973 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4199
  signal tmp_ivl_25974 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4199
  signal tmp_ivl_25979 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4199
  signal tmp_ivl_25981 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4199
  signal tmp_ivl_25986 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4200
  signal tmp_ivl_25991 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4200
  signal tmp_ivl_25993 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4200
  signal tmp_ivl_25998 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4200
  signal tmp_ivl_26000 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4200
  signal tmp_ivl_26005 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4201
  signal tmp_ivl_2601 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3029
  signal tmp_ivl_26010 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4201
  signal tmp_ivl_26013 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4201
  signal tmp_ivl_26014 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4201
  signal tmp_ivl_26019 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4201
  signal tmp_ivl_26021 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4201
  signal tmp_ivl_26027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4202
  signal tmp_ivl_26028 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4202
  signal tmp_ivl_2603 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3029
  signal tmp_ivl_26033 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4202
  signal tmp_ivl_26036 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4202
  signal tmp_ivl_26038 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4202
  signal tmp_ivl_26039 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4202
  signal tmp_ivl_26044 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4202
  signal tmp_ivl_26046 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4202
  signal tmp_ivl_2605 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3029
  signal tmp_ivl_26051 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4203
  signal tmp_ivl_26056 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4203
  signal tmp_ivl_26058 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4203
  signal tmp_ivl_26063 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4203
  signal tmp_ivl_26065 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4203
  signal tmp_ivl_26070 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4204
  signal tmp_ivl_26075 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4204
  signal tmp_ivl_26078 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4204
  signal tmp_ivl_26079 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4204
  signal tmp_ivl_26084 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4204
  signal tmp_ivl_26086 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4204
  signal tmp_ivl_26092 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4205
  signal tmp_ivl_26093 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4205
  signal tmp_ivl_26098 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4205
  signal tmp_ivl_26101 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4205
  signal tmp_ivl_26103 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4205
  signal tmp_ivl_26104 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4205
  signal tmp_ivl_26109 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4205
  signal tmp_ivl_2611 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3030
  signal tmp_ivl_26111 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4205
  signal tmp_ivl_26116 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4206
  signal tmp_ivl_26121 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4206
  signal tmp_ivl_26123 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4206
  signal tmp_ivl_26128 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4206
  signal tmp_ivl_2613 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3030
  signal tmp_ivl_26130 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4206
  signal tmp_ivl_26135 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4207
  signal tmp_ivl_2614 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3030
  signal tmp_ivl_26140 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4207
  signal tmp_ivl_26142 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4207
  signal tmp_ivl_26147 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4207
  signal tmp_ivl_26149 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4207
  signal tmp_ivl_26154 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4208
  signal tmp_ivl_26159 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4208
  signal tmp_ivl_26161 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4208
  signal tmp_ivl_26166 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4208
  signal tmp_ivl_26168 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4208
  signal tmp_ivl_26170 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4208
  signal tmp_ivl_26172 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4208
  signal tmp_ivl_26177 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4209
  signal tmp_ivl_26182 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4209
  signal tmp_ivl_26185 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4209
  signal tmp_ivl_26186 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4209
  signal tmp_ivl_2619 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3030
  signal tmp_ivl_26191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4209
  signal tmp_ivl_26193 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4209
  signal tmp_ivl_26199 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4210
  signal tmp_ivl_262 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2949
  signal tmp_ivl_26200 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4210
  signal tmp_ivl_26205 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4210
  signal tmp_ivl_26208 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4210
  signal tmp_ivl_26210 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4210
  signal tmp_ivl_26211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4210
  signal tmp_ivl_26216 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4210
  signal tmp_ivl_26218 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4210
  signal tmp_ivl_2622 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3030
  signal tmp_ivl_26223 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4211
  signal tmp_ivl_26228 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4211
  signal tmp_ivl_26230 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4211
  signal tmp_ivl_26235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4211
  signal tmp_ivl_26237 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4211
  signal tmp_ivl_2624 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3030
  signal tmp_ivl_26242 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4212
  signal tmp_ivl_26247 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4212
  signal tmp_ivl_2625 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3030
  signal tmp_ivl_26250 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4212
  signal tmp_ivl_26251 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4212
  signal tmp_ivl_26256 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4212
  signal tmp_ivl_26258 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4212
  signal tmp_ivl_26264 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4213
  signal tmp_ivl_26265 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4213
  signal tmp_ivl_26270 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4213
  signal tmp_ivl_26273 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4213
  signal tmp_ivl_26275 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4213
  signal tmp_ivl_26276 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4213
  signal tmp_ivl_26281 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4213
  signal tmp_ivl_26283 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4213
  signal tmp_ivl_26288 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4214
  signal tmp_ivl_26293 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4214
  signal tmp_ivl_26295 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4214
  signal tmp_ivl_2630 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3030
  signal tmp_ivl_26300 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4214
  signal tmp_ivl_26302 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4214
  signal tmp_ivl_26307 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4215
  signal tmp_ivl_26312 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4215
  signal tmp_ivl_26315 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4215
  signal tmp_ivl_26316 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4215
  signal tmp_ivl_2632 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3030
  signal tmp_ivl_26321 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4215
  signal tmp_ivl_26323 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4215
  signal tmp_ivl_26329 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4216
  signal tmp_ivl_26330 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4216
  signal tmp_ivl_26335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4216
  signal tmp_ivl_26338 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4216
  signal tmp_ivl_2634 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3030
  signal tmp_ivl_26340 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4216
  signal tmp_ivl_26341 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4216
  signal tmp_ivl_26346 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4216
  signal tmp_ivl_26348 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4216
  signal tmp_ivl_26353 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4217
  signal tmp_ivl_26358 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4217
  signal tmp_ivl_26360 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4217
  signal tmp_ivl_26365 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4217
  signal tmp_ivl_26367 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4217
  signal tmp_ivl_26372 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4218
  signal tmp_ivl_26377 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4218
  signal tmp_ivl_26379 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4218
  signal tmp_ivl_26384 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4218
  signal tmp_ivl_26386 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4218
  signal tmp_ivl_26391 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4219
  signal tmp_ivl_26396 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4219
  signal tmp_ivl_26398 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4219
  signal tmp_ivl_264 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2949
  signal tmp_ivl_2640 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3031
  signal tmp_ivl_26403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4219
  signal tmp_ivl_26405 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4219
  signal tmp_ivl_26407 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4219
  signal tmp_ivl_26409 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4219
  signal tmp_ivl_26414 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4220
  signal tmp_ivl_26419 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4220
  signal tmp_ivl_2642 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3031
  signal tmp_ivl_26422 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4220
  signal tmp_ivl_26423 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4220
  signal tmp_ivl_26428 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4220
  signal tmp_ivl_2643 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3031
  signal tmp_ivl_26430 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4220
  signal tmp_ivl_26436 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4221
  signal tmp_ivl_26437 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4221
  signal tmp_ivl_26442 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4221
  signal tmp_ivl_26445 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4221
  signal tmp_ivl_26447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4221
  signal tmp_ivl_26448 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4221
  signal tmp_ivl_26453 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4221
  signal tmp_ivl_26455 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4221
  signal tmp_ivl_26460 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4222
  signal tmp_ivl_26465 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4222
  signal tmp_ivl_26467 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4222
  signal tmp_ivl_26472 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4222
  signal tmp_ivl_26474 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4222
  signal tmp_ivl_26479 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4223
  signal tmp_ivl_2648 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3031
  signal tmp_ivl_26484 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4223
  signal tmp_ivl_26487 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4223
  signal tmp_ivl_26488 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4223
  signal tmp_ivl_26493 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4223
  signal tmp_ivl_26495 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4223
  signal tmp_ivl_265 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2949
  signal tmp_ivl_26501 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4224
  signal tmp_ivl_26502 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4224
  signal tmp_ivl_26507 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4224
  signal tmp_ivl_2651 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3031
  signal tmp_ivl_26510 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4224
  signal tmp_ivl_26512 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4224
  signal tmp_ivl_26513 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4224
  signal tmp_ivl_26518 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4224
  signal tmp_ivl_26520 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4224
  signal tmp_ivl_26525 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4225
  signal tmp_ivl_2653 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3031
  signal tmp_ivl_26530 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4225
  signal tmp_ivl_26532 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4225
  signal tmp_ivl_26537 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4225
  signal tmp_ivl_26539 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4225
  signal tmp_ivl_2654 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3031
  signal tmp_ivl_26544 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4226
  signal tmp_ivl_26549 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4226
  signal tmp_ivl_26551 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4226
  signal tmp_ivl_26556 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4226
  signal tmp_ivl_26558 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4226
  signal tmp_ivl_26563 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4227
  signal tmp_ivl_26568 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4227
  signal tmp_ivl_26571 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4227
  signal tmp_ivl_26572 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4227
  signal tmp_ivl_26577 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4227
  signal tmp_ivl_26579 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4227
  signal tmp_ivl_26585 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4228
  signal tmp_ivl_26586 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4228
  signal tmp_ivl_2659 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3031
  signal tmp_ivl_26591 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4228
  signal tmp_ivl_26594 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4228
  signal tmp_ivl_26596 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4228
  signal tmp_ivl_26597 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4228
  signal tmp_ivl_26602 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4228
  signal tmp_ivl_26604 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4228
  signal tmp_ivl_26609 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4229
  signal tmp_ivl_2661 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3031
  signal tmp_ivl_26614 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4229
  signal tmp_ivl_26616 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4229
  signal tmp_ivl_26621 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4229
  signal tmp_ivl_26623 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4229
  signal tmp_ivl_26628 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4230
  signal tmp_ivl_2663 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3031
  signal tmp_ivl_26633 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4230
  signal tmp_ivl_26635 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4230
  signal tmp_ivl_26640 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4230
  signal tmp_ivl_26642 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4230
  signal tmp_ivl_26644 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4230
  signal tmp_ivl_26646 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4230
  signal tmp_ivl_26651 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4231
  signal tmp_ivl_26656 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4231
  signal tmp_ivl_26659 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4231
  signal tmp_ivl_26660 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4231
  signal tmp_ivl_26665 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4231
  signal tmp_ivl_26667 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4231
  signal tmp_ivl_26673 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4232
  signal tmp_ivl_26674 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4232
  signal tmp_ivl_26679 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4232
  signal tmp_ivl_26682 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4232
  signal tmp_ivl_26684 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4232
  signal tmp_ivl_26685 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4232
  signal tmp_ivl_2669 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3032
  signal tmp_ivl_26690 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4232
  signal tmp_ivl_26692 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4232
  signal tmp_ivl_26697 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4233
  signal tmp_ivl_26702 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4233
  signal tmp_ivl_26704 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4233
  signal tmp_ivl_26709 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4233
  signal tmp_ivl_2671 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3032
  signal tmp_ivl_26711 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4233
  signal tmp_ivl_26716 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4234
  signal tmp_ivl_2672 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3032
  signal tmp_ivl_26721 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4234
  signal tmp_ivl_26724 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4234
  signal tmp_ivl_26725 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4234
  signal tmp_ivl_26730 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4234
  signal tmp_ivl_26732 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4234
  signal tmp_ivl_26738 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4235
  signal tmp_ivl_26739 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4235
  signal tmp_ivl_26744 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4235
  signal tmp_ivl_26747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4235
  signal tmp_ivl_26749 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4235
  signal tmp_ivl_26750 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4235
  signal tmp_ivl_26755 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4235
  signal tmp_ivl_26757 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4235
  signal tmp_ivl_26762 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4236
  signal tmp_ivl_26767 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4236
  signal tmp_ivl_26769 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4236
  signal tmp_ivl_2677 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3032
  signal tmp_ivl_26774 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4236
  signal tmp_ivl_26776 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4236
  signal tmp_ivl_26781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4237
  signal tmp_ivl_26786 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4237
  signal tmp_ivl_26788 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4237
  signal tmp_ivl_26793 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4237
  signal tmp_ivl_26795 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4237
  signal tmp_ivl_2680 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3032
  signal tmp_ivl_26800 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4238
  signal tmp_ivl_26805 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4238
  signal tmp_ivl_26808 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4238
  signal tmp_ivl_26809 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4238
  signal tmp_ivl_26814 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4238
  signal tmp_ivl_26816 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4238
  signal tmp_ivl_2682 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3032
  signal tmp_ivl_26822 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4239
  signal tmp_ivl_26823 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4239
  signal tmp_ivl_26828 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4239
  signal tmp_ivl_2683 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3032
  signal tmp_ivl_26831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4239
  signal tmp_ivl_26833 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4239
  signal tmp_ivl_26834 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4239
  signal tmp_ivl_26839 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4239
  signal tmp_ivl_26841 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4239
  signal tmp_ivl_26846 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4240
  signal tmp_ivl_26851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4240
  signal tmp_ivl_26853 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4240
  signal tmp_ivl_26858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4240
  signal tmp_ivl_26860 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4240
  signal tmp_ivl_26865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4241
  signal tmp_ivl_26870 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4241
  signal tmp_ivl_26872 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4241
  signal tmp_ivl_26877 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4241
  signal tmp_ivl_26879 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4241
  signal tmp_ivl_2688 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3032
  signal tmp_ivl_26881 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4241
  signal tmp_ivl_26883 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4241
  signal tmp_ivl_26888 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4242
  signal tmp_ivl_26893 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4242
  signal tmp_ivl_26896 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4242
  signal tmp_ivl_26897 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4242
  signal tmp_ivl_2690 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3032
  signal tmp_ivl_26902 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4242
  signal tmp_ivl_26904 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4242
  signal tmp_ivl_26910 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4243
  signal tmp_ivl_26911 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4243
  signal tmp_ivl_26916 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4243
  signal tmp_ivl_26919 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4243
  signal tmp_ivl_2692 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3032
  signal tmp_ivl_26921 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4243
  signal tmp_ivl_26922 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4243
  signal tmp_ivl_26927 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4243
  signal tmp_ivl_26929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4243
  signal tmp_ivl_26934 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4244
  signal tmp_ivl_26939 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4244
  signal tmp_ivl_26941 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4244
  signal tmp_ivl_26946 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4244
  signal tmp_ivl_26948 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4244
  signal tmp_ivl_26953 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4245
  signal tmp_ivl_26958 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4245
  signal tmp_ivl_26961 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4245
  signal tmp_ivl_26962 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4245
  signal tmp_ivl_26967 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4245
  signal tmp_ivl_26969 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4245
  signal tmp_ivl_26975 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4246
  signal tmp_ivl_26976 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4246
  signal tmp_ivl_2698 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3033
  signal tmp_ivl_26981 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4246
  signal tmp_ivl_26984 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4246
  signal tmp_ivl_26986 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4246
  signal tmp_ivl_26987 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4246
  signal tmp_ivl_26992 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4246
  signal tmp_ivl_26994 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4246
  signal tmp_ivl_26999 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4247
  signal tmp_ivl_270 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2949
  signal tmp_ivl_2700 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3033
  signal tmp_ivl_27004 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4247
  signal tmp_ivl_27006 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4247
  signal tmp_ivl_2701 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3033
  signal tmp_ivl_27011 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4247
  signal tmp_ivl_27013 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4247
  signal tmp_ivl_27018 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4248
  signal tmp_ivl_27023 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4248
  signal tmp_ivl_27026 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4248
  signal tmp_ivl_27027 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4248
  signal tmp_ivl_27032 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4248
  signal tmp_ivl_27034 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4248
  signal tmp_ivl_27040 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4249
  signal tmp_ivl_27041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4249
  signal tmp_ivl_27046 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4249
  signal tmp_ivl_27049 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4249
  signal tmp_ivl_27051 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4249
  signal tmp_ivl_27052 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4249
  signal tmp_ivl_27057 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4249
  signal tmp_ivl_27059 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4249
  signal tmp_ivl_2706 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3033
  signal tmp_ivl_27064 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4250
  signal tmp_ivl_27069 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4250
  signal tmp_ivl_27071 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4250
  signal tmp_ivl_27076 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4250
  signal tmp_ivl_27078 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4250
  signal tmp_ivl_27083 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4251
  signal tmp_ivl_27088 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4251
  signal tmp_ivl_2709 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3033
  signal tmp_ivl_27090 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4251
  signal tmp_ivl_27095 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4251
  signal tmp_ivl_27097 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4251
  signal tmp_ivl_27102 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4252
  signal tmp_ivl_27107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4252
  signal tmp_ivl_27109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4252
  signal tmp_ivl_2711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3033
  signal tmp_ivl_27114 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4252
  signal tmp_ivl_27116 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4252
  signal tmp_ivl_27118 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4252
  signal tmp_ivl_2712 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3033
  signal tmp_ivl_27120 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4252
  signal tmp_ivl_27125 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4253
  signal tmp_ivl_27130 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4253
  signal tmp_ivl_27133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4253
  signal tmp_ivl_27134 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4253
  signal tmp_ivl_27139 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4253
  signal tmp_ivl_27141 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4253
  signal tmp_ivl_27147 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4254
  signal tmp_ivl_27148 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4254
  signal tmp_ivl_27153 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4254
  signal tmp_ivl_27156 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4254
  signal tmp_ivl_27158 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4254
  signal tmp_ivl_27159 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4254
  signal tmp_ivl_27164 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4254
  signal tmp_ivl_27166 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4254
  signal tmp_ivl_2717 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3033
  signal tmp_ivl_27171 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4255
  signal tmp_ivl_27176 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4255
  signal tmp_ivl_27178 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4255
  signal tmp_ivl_27183 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4255
  signal tmp_ivl_27185 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4255
  signal tmp_ivl_2719 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3033
  signal tmp_ivl_27190 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4256
  signal tmp_ivl_27195 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4256
  signal tmp_ivl_27197 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4256
  signal tmp_ivl_27202 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4256
  signal tmp_ivl_27204 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4256
  signal tmp_ivl_27209 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4257
  signal tmp_ivl_2721 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3033
  signal tmp_ivl_27214 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4257
  signal tmp_ivl_27217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4257
  signal tmp_ivl_27218 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4257
  signal tmp_ivl_27223 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4257
  signal tmp_ivl_27225 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4257
  signal tmp_ivl_27231 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4258
  signal tmp_ivl_27232 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4258
  signal tmp_ivl_27237 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4258
  signal tmp_ivl_27240 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4258
  signal tmp_ivl_27242 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4258
  signal tmp_ivl_27243 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4258
  signal tmp_ivl_27248 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4258
  signal tmp_ivl_27250 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4258
  signal tmp_ivl_27255 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4259
  signal tmp_ivl_27260 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4259
  signal tmp_ivl_27262 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4259
  signal tmp_ivl_27267 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4259
  signal tmp_ivl_27269 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4259
  signal tmp_ivl_2727 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3034
  signal tmp_ivl_27274 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4260
  signal tmp_ivl_27279 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4260
  signal tmp_ivl_27281 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4260
  signal tmp_ivl_27286 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4260
  signal tmp_ivl_27288 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4260
  signal tmp_ivl_2729 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3034
  signal tmp_ivl_27290 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4260
  signal tmp_ivl_27292 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4260
  signal tmp_ivl_27297 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4261
  signal tmp_ivl_273 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2949
  signal tmp_ivl_2730 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3034
  signal tmp_ivl_27302 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4261
  signal tmp_ivl_27305 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4261
  signal tmp_ivl_27306 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4261
  signal tmp_ivl_27311 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4261
  signal tmp_ivl_27313 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4261
  signal tmp_ivl_27319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4262
  signal tmp_ivl_27320 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4262
  signal tmp_ivl_27325 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4262
  signal tmp_ivl_27328 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4262
  signal tmp_ivl_27330 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4262
  signal tmp_ivl_27331 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4262
  signal tmp_ivl_27336 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4262
  signal tmp_ivl_27338 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4262
  signal tmp_ivl_27343 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4263
  signal tmp_ivl_27348 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4263
  signal tmp_ivl_2735 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3034
  signal tmp_ivl_27350 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4263
  signal tmp_ivl_27355 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4263
  signal tmp_ivl_27357 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4263
  signal tmp_ivl_27362 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4264
  signal tmp_ivl_27367 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4264
  signal tmp_ivl_27369 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4264
  signal tmp_ivl_27374 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4264
  signal tmp_ivl_27376 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4264
  signal tmp_ivl_2738 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3034
  signal tmp_ivl_27381 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4265
  signal tmp_ivl_27386 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4265
  signal tmp_ivl_27389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4265
  signal tmp_ivl_27390 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4265
  signal tmp_ivl_27395 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4265
  signal tmp_ivl_27397 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4265
  signal tmp_ivl_2740 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3034
  signal tmp_ivl_27403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4266
  signal tmp_ivl_27404 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4266
  signal tmp_ivl_27409 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4266
  signal tmp_ivl_2741 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3034
  signal tmp_ivl_27412 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4266
  signal tmp_ivl_27414 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4266
  signal tmp_ivl_27415 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4266
  signal tmp_ivl_27420 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4266
  signal tmp_ivl_27422 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4266
  signal tmp_ivl_27427 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4267
  signal tmp_ivl_27432 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4267
  signal tmp_ivl_27434 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4267
  signal tmp_ivl_27439 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4267
  signal tmp_ivl_27441 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4267
  signal tmp_ivl_27446 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4268
  signal tmp_ivl_27451 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4268
  signal tmp_ivl_27453 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4268
  signal tmp_ivl_27458 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4268
  signal tmp_ivl_2746 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3034
  signal tmp_ivl_27460 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4268
  signal tmp_ivl_27462 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4268
  signal tmp_ivl_27464 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4268
  signal tmp_ivl_27469 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4269
  signal tmp_ivl_27474 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4269
  signal tmp_ivl_27477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4269
  signal tmp_ivl_27478 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4269
  signal tmp_ivl_2748 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3034
  signal tmp_ivl_27483 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4269
  signal tmp_ivl_27485 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4269
  signal tmp_ivl_27491 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4270
  signal tmp_ivl_27492 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4270
  signal tmp_ivl_27497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4270
  signal tmp_ivl_275 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2949
  signal tmp_ivl_2750 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3034
  signal tmp_ivl_27500 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4270
  signal tmp_ivl_27502 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4270
  signal tmp_ivl_27503 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4270
  signal tmp_ivl_27508 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4270
  signal tmp_ivl_27510 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4270
  signal tmp_ivl_27515 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4271
  signal tmp_ivl_27520 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4271
  signal tmp_ivl_27522 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4271
  signal tmp_ivl_27527 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4271
  signal tmp_ivl_27529 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4271
  signal tmp_ivl_27534 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4272
  signal tmp_ivl_27539 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4272
  signal tmp_ivl_27542 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4272
  signal tmp_ivl_27543 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4272
  signal tmp_ivl_27548 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4272
  signal tmp_ivl_27550 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4272
  signal tmp_ivl_27556 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4273
  signal tmp_ivl_27557 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4273
  signal tmp_ivl_2756 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3035
  signal tmp_ivl_27562 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4273
  signal tmp_ivl_27565 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4273
  signal tmp_ivl_27567 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4273
  signal tmp_ivl_27568 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4273
  signal tmp_ivl_27573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4273
  signal tmp_ivl_27575 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4273
  signal tmp_ivl_2758 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3035
  signal tmp_ivl_27580 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4274
  signal tmp_ivl_27585 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4274
  signal tmp_ivl_27587 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4274
  signal tmp_ivl_2759 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3035
  signal tmp_ivl_27592 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4274
  signal tmp_ivl_27594 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4274
  signal tmp_ivl_27599 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4275
  signal tmp_ivl_276 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2949
  signal tmp_ivl_27604 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4275
  signal tmp_ivl_27606 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4275
  signal tmp_ivl_27611 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4275
  signal tmp_ivl_27613 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4275
  signal tmp_ivl_27618 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4276
  signal tmp_ivl_27623 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4276
  signal tmp_ivl_27625 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4276
  signal tmp_ivl_27630 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4276
  signal tmp_ivl_27632 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4276
  signal tmp_ivl_27634 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4276
  signal tmp_ivl_27636 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4276
  signal tmp_ivl_2764 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3035
  signal tmp_ivl_27641 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4277
  signal tmp_ivl_27646 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4277
  signal tmp_ivl_27648 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4277
  signal tmp_ivl_27653 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4277
  signal tmp_ivl_27655 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4277
  signal tmp_ivl_27660 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4278
  signal tmp_ivl_27665 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4278
  signal tmp_ivl_27668 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4278
  signal tmp_ivl_27669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4278
  signal tmp_ivl_2767 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3035
  signal tmp_ivl_27674 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4278
  signal tmp_ivl_27676 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4278
  signal tmp_ivl_27682 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4279
  signal tmp_ivl_27683 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4279
  signal tmp_ivl_27688 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4279
  signal tmp_ivl_2769 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3035
  signal tmp_ivl_27691 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4279
  signal tmp_ivl_27693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4279
  signal tmp_ivl_27694 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4279
  signal tmp_ivl_27699 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4279
  signal tmp_ivl_2770 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3035
  signal tmp_ivl_27701 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4279
  signal tmp_ivl_27706 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4280
  signal tmp_ivl_27711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4280
  signal tmp_ivl_27713 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4280
  signal tmp_ivl_27718 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4280
  signal tmp_ivl_27720 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4280
  signal tmp_ivl_27725 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4281
  signal tmp_ivl_27730 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4281
  signal tmp_ivl_27732 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4281
  signal tmp_ivl_27737 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4281
  signal tmp_ivl_27739 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4281
  signal tmp_ivl_27741 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4281
  signal tmp_ivl_27743 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4281
  signal tmp_ivl_27748 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4282
  signal tmp_ivl_2775 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3035
  signal tmp_ivl_27753 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4282
  signal tmp_ivl_27755 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4282
  signal tmp_ivl_27760 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4282
  signal tmp_ivl_27762 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4282
  signal tmp_ivl_27767 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4283
  signal tmp_ivl_2777 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3035
  signal tmp_ivl_27772 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4283
  signal tmp_ivl_27775 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4283
  signal tmp_ivl_27776 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4283
  signal tmp_ivl_27781 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4283
  signal tmp_ivl_27783 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4283
  signal tmp_ivl_27789 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4284
  signal tmp_ivl_2779 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3035
  signal tmp_ivl_27790 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4284
  signal tmp_ivl_27795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4284
  signal tmp_ivl_27798 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4284
  signal tmp_ivl_27800 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4284
  signal tmp_ivl_27801 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4284
  signal tmp_ivl_27806 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4284
  signal tmp_ivl_27808 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4284
  signal tmp_ivl_27813 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4285
  signal tmp_ivl_27818 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4285
  signal tmp_ivl_27820 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4285
  signal tmp_ivl_27825 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4285
  signal tmp_ivl_27827 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4285
  signal tmp_ivl_27832 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4286
  signal tmp_ivl_27837 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4286
  signal tmp_ivl_27839 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4286
  signal tmp_ivl_27844 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4286
  signal tmp_ivl_27846 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4286
  signal tmp_ivl_27848 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4286
  signal tmp_ivl_2785 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3036
  signal tmp_ivl_27850 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4286
  signal tmp_ivl_27855 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4287
  signal tmp_ivl_27860 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4287
  signal tmp_ivl_27862 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4287
  signal tmp_ivl_27867 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4287
  signal tmp_ivl_27869 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4287
  signal tmp_ivl_2787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3036
  signal tmp_ivl_27874 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4288
  signal tmp_ivl_27879 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4288
  signal tmp_ivl_2788 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3036
  signal tmp_ivl_27882 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4288
  signal tmp_ivl_27883 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4288
  signal tmp_ivl_27888 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4288
  signal tmp_ivl_27890 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4288
  signal tmp_ivl_27896 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4289
  signal tmp_ivl_27897 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4289
  signal tmp_ivl_27902 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4289
  signal tmp_ivl_27905 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4289
  signal tmp_ivl_27907 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4289
  signal tmp_ivl_27908 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4289
  signal tmp_ivl_27913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4289
  signal tmp_ivl_27915 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4289
  signal tmp_ivl_27920 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4290
  signal tmp_ivl_27925 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4290
  signal tmp_ivl_27927 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4290
  signal tmp_ivl_2793 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3036
  signal tmp_ivl_27932 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4290
  signal tmp_ivl_27934 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4290
  signal tmp_ivl_27939 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4291
  signal tmp_ivl_27944 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4291
  signal tmp_ivl_27946 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4291
  signal tmp_ivl_27951 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4291
  signal tmp_ivl_27953 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4291
  signal tmp_ivl_27955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4291
  signal tmp_ivl_27957 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4291
  signal tmp_ivl_2796 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3036
  signal tmp_ivl_27962 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4292
  signal tmp_ivl_27967 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4292
  signal tmp_ivl_27969 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4292
  signal tmp_ivl_27974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4292
  signal tmp_ivl_27976 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4292
  signal tmp_ivl_2798 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3036
  signal tmp_ivl_27981 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4293
  signal tmp_ivl_27986 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4293
  signal tmp_ivl_27989 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4293
  signal tmp_ivl_2799 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3036
  signal tmp_ivl_27990 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4293
  signal tmp_ivl_27995 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4293
  signal tmp_ivl_27997 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4293
  signal tmp_ivl_28003 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4294
  signal tmp_ivl_28004 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4294
  signal tmp_ivl_28009 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4294
  signal tmp_ivl_28012 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4294
  signal tmp_ivl_28014 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4294
  signal tmp_ivl_28015 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4294
  signal tmp_ivl_28020 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4294
  signal tmp_ivl_28022 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4294
  signal tmp_ivl_28027 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4295
  signal tmp_ivl_28032 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4295
  signal tmp_ivl_28034 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4295
  signal tmp_ivl_28039 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4295
  signal tmp_ivl_2804 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3036
  signal tmp_ivl_28041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4295
  signal tmp_ivl_28046 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4296
  signal tmp_ivl_28051 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4296
  signal tmp_ivl_28053 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4296
  signal tmp_ivl_28058 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4296
  signal tmp_ivl_2806 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3036
  signal tmp_ivl_28060 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4296
  signal tmp_ivl_28062 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4296
  signal tmp_ivl_28064 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4296
  signal tmp_ivl_28069 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4297
  signal tmp_ivl_28074 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4297
  signal tmp_ivl_28076 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4297
  signal tmp_ivl_2808 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3036
  signal tmp_ivl_28081 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4297
  signal tmp_ivl_28083 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4297
  signal tmp_ivl_28088 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4298
  signal tmp_ivl_28093 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4298
  signal tmp_ivl_28096 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4298
  signal tmp_ivl_28097 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4298
  signal tmp_ivl_281 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2949
  signal tmp_ivl_28102 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4298
  signal tmp_ivl_28104 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4298
  signal tmp_ivl_28110 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4299
  signal tmp_ivl_28111 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4299
  signal tmp_ivl_28116 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4299
  signal tmp_ivl_28119 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4299
  signal tmp_ivl_28121 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4299
  signal tmp_ivl_28122 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4299
  signal tmp_ivl_28127 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4299
  signal tmp_ivl_28129 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4299
  signal tmp_ivl_28134 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4300
  signal tmp_ivl_28139 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4300
  signal tmp_ivl_2814 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3037
  signal tmp_ivl_28141 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4300
  signal tmp_ivl_28146 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4300
  signal tmp_ivl_28148 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4300
  signal tmp_ivl_28153 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4301
  signal tmp_ivl_28158 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4301
  signal tmp_ivl_2816 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3037
  signal tmp_ivl_28160 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4301
  signal tmp_ivl_28165 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4301
  signal tmp_ivl_28167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4301
  signal tmp_ivl_28169 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4301
  signal tmp_ivl_2817 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3037
  signal tmp_ivl_28171 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4301
  signal tmp_ivl_28176 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4302
  signal tmp_ivl_28181 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4302
  signal tmp_ivl_28183 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4302
  signal tmp_ivl_28188 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4302
  signal tmp_ivl_28190 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4302
  signal tmp_ivl_28195 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4303
  signal tmp_ivl_28200 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4303
  signal tmp_ivl_28203 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4303
  signal tmp_ivl_28204 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4303
  signal tmp_ivl_28209 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4303
  signal tmp_ivl_28211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4303
  signal tmp_ivl_28217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4304
  signal tmp_ivl_28218 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4304
  signal tmp_ivl_2822 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3037
  signal tmp_ivl_28223 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4304
  signal tmp_ivl_28226 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4304
  signal tmp_ivl_28228 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4304
  signal tmp_ivl_28229 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4304
  signal tmp_ivl_28234 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4304
  signal tmp_ivl_28236 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4304
  signal tmp_ivl_28241 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4305
  signal tmp_ivl_28246 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4305
  signal tmp_ivl_28248 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4305
  signal tmp_ivl_2825 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3037
  signal tmp_ivl_28253 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4305
  signal tmp_ivl_28255 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4305
  signal tmp_ivl_28260 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4306
  signal tmp_ivl_28265 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4306
  signal tmp_ivl_28267 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4306
  signal tmp_ivl_2827 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3037
  signal tmp_ivl_28272 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4306
  signal tmp_ivl_28274 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4306
  signal tmp_ivl_28276 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4306
  signal tmp_ivl_28278 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4306
  signal tmp_ivl_2828 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3037
  signal tmp_ivl_28283 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4307
  signal tmp_ivl_28288 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4307
  signal tmp_ivl_28290 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4307
  signal tmp_ivl_28295 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4307
  signal tmp_ivl_28297 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4307
  signal tmp_ivl_283 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2949
  signal tmp_ivl_28302 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4308
  signal tmp_ivl_28307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4308
  signal tmp_ivl_28310 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4308
  signal tmp_ivl_28311 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4308
  signal tmp_ivl_28316 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4308
  signal tmp_ivl_28318 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4308
  signal tmp_ivl_28324 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4309
  signal tmp_ivl_28325 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4309
  signal tmp_ivl_2833 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3037
  signal tmp_ivl_28330 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4309
  signal tmp_ivl_28333 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4309
  signal tmp_ivl_28335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4309
  signal tmp_ivl_28336 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4309
  signal tmp_ivl_28341 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4309
  signal tmp_ivl_28343 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4309
  signal tmp_ivl_28348 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4310
  signal tmp_ivl_2835 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3037
  signal tmp_ivl_28353 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4310
  signal tmp_ivl_28355 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4310
  signal tmp_ivl_28360 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4310
  signal tmp_ivl_28362 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4310
  signal tmp_ivl_28367 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4311
  signal tmp_ivl_2837 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3037
  signal tmp_ivl_28372 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4311
  signal tmp_ivl_28374 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4311
  signal tmp_ivl_28379 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4311
  signal tmp_ivl_28381 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4311
  signal tmp_ivl_28383 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4311
  signal tmp_ivl_28385 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4311
  signal tmp_ivl_28390 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4312
  signal tmp_ivl_28395 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4312
  signal tmp_ivl_28398 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4312
  signal tmp_ivl_28399 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4312
  signal tmp_ivl_28404 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4312
  signal tmp_ivl_28406 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4312
  signal tmp_ivl_28412 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4313
  signal tmp_ivl_28413 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4313
  signal tmp_ivl_28418 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4313
  signal tmp_ivl_28421 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4313
  signal tmp_ivl_28423 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4313
  signal tmp_ivl_28424 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4313
  signal tmp_ivl_28429 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4313
  signal tmp_ivl_2843 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3038
  signal tmp_ivl_28431 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4313
  signal tmp_ivl_28436 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4314
  signal tmp_ivl_28441 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4314
  signal tmp_ivl_28443 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4314
  signal tmp_ivl_28448 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4314
  signal tmp_ivl_2845 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3038
  signal tmp_ivl_28450 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4314
  signal tmp_ivl_28455 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4315
  signal tmp_ivl_2846 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3038
  signal tmp_ivl_28460 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4315
  signal tmp_ivl_28462 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4315
  signal tmp_ivl_28467 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4315
  signal tmp_ivl_28469 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4315
  signal tmp_ivl_28474 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4316
  signal tmp_ivl_28479 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4316
  signal tmp_ivl_28481 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4316
  signal tmp_ivl_28486 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4316
  signal tmp_ivl_28488 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4316
  signal tmp_ivl_28490 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4316
  signal tmp_ivl_28492 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4316
  signal tmp_ivl_28497 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4317
  signal tmp_ivl_285 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2949
  signal tmp_ivl_28502 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4317
  signal tmp_ivl_28505 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4317
  signal tmp_ivl_28506 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4317
  signal tmp_ivl_2851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3038
  signal tmp_ivl_28511 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4317
  signal tmp_ivl_28513 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4317
  signal tmp_ivl_28519 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4318
  signal tmp_ivl_28520 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4318
  signal tmp_ivl_28525 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4318
  signal tmp_ivl_28528 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4318
  signal tmp_ivl_28530 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4318
  signal tmp_ivl_28531 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4318
  signal tmp_ivl_28536 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4318
  signal tmp_ivl_28538 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4318
  signal tmp_ivl_2854 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3038
  signal tmp_ivl_28543 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4319
  signal tmp_ivl_28548 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4319
  signal tmp_ivl_28550 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4319
  signal tmp_ivl_28555 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4319
  signal tmp_ivl_28557 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4319
  signal tmp_ivl_2856 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3038
  signal tmp_ivl_28562 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4320
  signal tmp_ivl_28567 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4320
  signal tmp_ivl_28569 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4320
  signal tmp_ivl_2857 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3038
  signal tmp_ivl_28574 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4320
  signal tmp_ivl_28576 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4320
  signal tmp_ivl_28581 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4321
  signal tmp_ivl_28586 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4321
  signal tmp_ivl_28588 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4321
  signal tmp_ivl_28593 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4321
  signal tmp_ivl_28595 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4321
  signal tmp_ivl_28597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4321
  signal tmp_ivl_28599 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4321
  signal tmp_ivl_28604 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4322
  signal tmp_ivl_28609 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4322
  signal tmp_ivl_28611 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4322
  signal tmp_ivl_28616 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4322
  signal tmp_ivl_28618 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4322
  signal tmp_ivl_2862 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3038
  signal tmp_ivl_28623 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4323
  signal tmp_ivl_28628 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4323
  signal tmp_ivl_28631 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4323
  signal tmp_ivl_28632 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4323
  signal tmp_ivl_28637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4323
  signal tmp_ivl_28639 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4323
  signal tmp_ivl_2864 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3038
  signal tmp_ivl_28645 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4324
  signal tmp_ivl_28646 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4324
  signal tmp_ivl_28651 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4324
  signal tmp_ivl_28654 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4324
  signal tmp_ivl_28656 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4324
  signal tmp_ivl_28657 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4324
  signal tmp_ivl_2866 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3038
  signal tmp_ivl_28662 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4324
  signal tmp_ivl_28664 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4324
  signal tmp_ivl_28669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4325
  signal tmp_ivl_28674 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4325
  signal tmp_ivl_28676 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4325
  signal tmp_ivl_28681 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4325
  signal tmp_ivl_28683 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4325
  signal tmp_ivl_28688 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4326
  signal tmp_ivl_28693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4326
  signal tmp_ivl_28695 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4326
  signal tmp_ivl_28700 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4326
  signal tmp_ivl_28702 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4326
  signal tmp_ivl_28704 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4326
  signal tmp_ivl_28706 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4326
  signal tmp_ivl_28711 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4327
  signal tmp_ivl_28716 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4327
  signal tmp_ivl_28718 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4327
  signal tmp_ivl_2872 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3039
  signal tmp_ivl_28723 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4327
  signal tmp_ivl_28725 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4327
  signal tmp_ivl_28730 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4328
  signal tmp_ivl_28735 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4328
  signal tmp_ivl_28738 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4328
  signal tmp_ivl_28739 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4328
  signal tmp_ivl_2874 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3039
  signal tmp_ivl_28744 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4328
  signal tmp_ivl_28746 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4328
  signal tmp_ivl_2875 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3039
  signal tmp_ivl_28752 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4329
  signal tmp_ivl_28753 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4329
  signal tmp_ivl_28758 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4329
  signal tmp_ivl_28761 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4329
  signal tmp_ivl_28763 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4329
  signal tmp_ivl_28764 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4329
  signal tmp_ivl_28769 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4329
  signal tmp_ivl_28771 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4329
  signal tmp_ivl_28776 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4330
  signal tmp_ivl_28781 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4330
  signal tmp_ivl_28783 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4330
  signal tmp_ivl_28788 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4330
  signal tmp_ivl_28790 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4330
  signal tmp_ivl_28795 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4331
  signal tmp_ivl_2880 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3039
  signal tmp_ivl_28800 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4331
  signal tmp_ivl_28802 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4331
  signal tmp_ivl_28807 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4331
  signal tmp_ivl_28809 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4331
  signal tmp_ivl_28811 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4331
  signal tmp_ivl_28813 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4331
  signal tmp_ivl_28818 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4332
  signal tmp_ivl_28823 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4332
  signal tmp_ivl_28826 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4332
  signal tmp_ivl_28827 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4332
  signal tmp_ivl_2883 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3039
  signal tmp_ivl_28832 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4332
  signal tmp_ivl_28834 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4332
  signal tmp_ivl_28840 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4333
  signal tmp_ivl_28841 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4333
  signal tmp_ivl_28846 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4333
  signal tmp_ivl_28849 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4333
  signal tmp_ivl_2885 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3039
  signal tmp_ivl_28851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4333
  signal tmp_ivl_28852 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4333
  signal tmp_ivl_28857 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4333
  signal tmp_ivl_28859 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4333
  signal tmp_ivl_2886 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3039
  signal tmp_ivl_28864 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4334
  signal tmp_ivl_28869 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4334
  signal tmp_ivl_28871 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4334
  signal tmp_ivl_28876 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4334
  signal tmp_ivl_28878 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4334
  signal tmp_ivl_28883 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4335
  signal tmp_ivl_28888 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4335
  signal tmp_ivl_28890 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4335
  signal tmp_ivl_28895 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4335
  signal tmp_ivl_28897 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4335
  signal tmp_ivl_28902 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4336
  signal tmp_ivl_28907 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4336
  signal tmp_ivl_28909 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4336
  signal tmp_ivl_2891 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3039
  signal tmp_ivl_28914 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4336
  signal tmp_ivl_28916 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4336
  signal tmp_ivl_28918 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4336
  signal tmp_ivl_28920 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4336
  signal tmp_ivl_28925 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4337
  signal tmp_ivl_2893 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3039
  signal tmp_ivl_28930 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4337
  signal tmp_ivl_28932 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4337
  signal tmp_ivl_28937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4337
  signal tmp_ivl_28939 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4337
  signal tmp_ivl_28944 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4338
  signal tmp_ivl_28949 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4338
  signal tmp_ivl_2895 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3039
  signal tmp_ivl_28952 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4338
  signal tmp_ivl_28953 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4338
  signal tmp_ivl_28958 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4338
  signal tmp_ivl_28960 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4338
  signal tmp_ivl_28966 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4339
  signal tmp_ivl_28967 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4339
  signal tmp_ivl_28972 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4339
  signal tmp_ivl_28975 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4339
  signal tmp_ivl_28977 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4339
  signal tmp_ivl_28978 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4339
  signal tmp_ivl_28983 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4339
  signal tmp_ivl_28985 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4339
  signal tmp_ivl_28990 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4340
  signal tmp_ivl_28995 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4340
  signal tmp_ivl_28997 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4340
  signal tmp_ivl_29002 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4340
  signal tmp_ivl_29004 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4340
  signal tmp_ivl_29009 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4341
  signal tmp_ivl_2901 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3040
  signal tmp_ivl_29014 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4341
  signal tmp_ivl_29016 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4341
  signal tmp_ivl_29021 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4341
  signal tmp_ivl_29023 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4341
  signal tmp_ivl_29025 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4341
  signal tmp_ivl_29027 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4341
  signal tmp_ivl_2903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3040
  signal tmp_ivl_29032 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4342
  signal tmp_ivl_29037 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4342
  signal tmp_ivl_2904 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3040
  signal tmp_ivl_29040 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4342
  signal tmp_ivl_29041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4342
  signal tmp_ivl_29046 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4342
  signal tmp_ivl_29048 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4342
  signal tmp_ivl_29054 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4343
  signal tmp_ivl_29055 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4343
  signal tmp_ivl_29060 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4343
  signal tmp_ivl_29063 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4343
  signal tmp_ivl_29065 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4343
  signal tmp_ivl_29066 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4343
  signal tmp_ivl_29071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4343
  signal tmp_ivl_29073 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4343
  signal tmp_ivl_29078 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4344
  signal tmp_ivl_29083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4344
  signal tmp_ivl_29085 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4344
  signal tmp_ivl_2909 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3040
  signal tmp_ivl_29090 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4344
  signal tmp_ivl_29092 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4344
  signal tmp_ivl_29097 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4345
  signal tmp_ivl_291 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2950
  signal tmp_ivl_29102 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4345
  signal tmp_ivl_29104 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4345
  signal tmp_ivl_29109 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4345
  signal tmp_ivl_29111 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4345
  signal tmp_ivl_29116 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4346
  signal tmp_ivl_2912 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3040
  signal tmp_ivl_29121 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4346
  signal tmp_ivl_29123 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4346
  signal tmp_ivl_29128 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4346
  signal tmp_ivl_29130 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4346
  signal tmp_ivl_29132 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4346
  signal tmp_ivl_29134 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4346
  signal tmp_ivl_29139 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4347
  signal tmp_ivl_2914 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3040
  signal tmp_ivl_29144 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4347
  signal tmp_ivl_29147 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4347
  signal tmp_ivl_29148 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4347
  signal tmp_ivl_2915 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3040
  signal tmp_ivl_29153 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4347
  signal tmp_ivl_29155 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4347
  signal tmp_ivl_29161 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4348
  signal tmp_ivl_29162 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4348
  signal tmp_ivl_29167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4348
  signal tmp_ivl_29170 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4348
  signal tmp_ivl_29172 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4348
  signal tmp_ivl_29173 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4348
  signal tmp_ivl_29178 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4348
  signal tmp_ivl_29180 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4348
  signal tmp_ivl_29185 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4349
  signal tmp_ivl_29190 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4349
  signal tmp_ivl_29192 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4349
  signal tmp_ivl_29197 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4349
  signal tmp_ivl_29199 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4349
  signal tmp_ivl_2920 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3040
  signal tmp_ivl_29204 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4350
  signal tmp_ivl_29209 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4350
  signal tmp_ivl_29211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4350
  signal tmp_ivl_29216 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4350
  signal tmp_ivl_29218 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4350
  signal tmp_ivl_2922 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3040
  signal tmp_ivl_29223 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4351
  signal tmp_ivl_29228 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4351
  signal tmp_ivl_29230 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4351
  signal tmp_ivl_29235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4351
  signal tmp_ivl_29237 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4351
  signal tmp_ivl_29239 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4351
  signal tmp_ivl_2924 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3040
  signal tmp_ivl_29241 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4351
  signal tmp_ivl_29246 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4352
  signal tmp_ivl_29251 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4352
  signal tmp_ivl_29253 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4352
  signal tmp_ivl_29258 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4352
  signal tmp_ivl_29260 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4352
  signal tmp_ivl_29265 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4353
  signal tmp_ivl_29270 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4353
  signal tmp_ivl_29273 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4353
  signal tmp_ivl_29274 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4353
  signal tmp_ivl_29279 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4353
  signal tmp_ivl_29281 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4353
  signal tmp_ivl_29287 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4354
  signal tmp_ivl_29288 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4354
  signal tmp_ivl_29293 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4354
  signal tmp_ivl_29296 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4354
  signal tmp_ivl_29298 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4354
  signal tmp_ivl_29299 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4354
  signal tmp_ivl_293 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2950
  signal tmp_ivl_2930 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3041
  signal tmp_ivl_29304 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4354
  signal tmp_ivl_29306 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4354
  signal tmp_ivl_29311 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4355
  signal tmp_ivl_29316 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4355
  signal tmp_ivl_29318 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4355
  signal tmp_ivl_2932 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3041
  signal tmp_ivl_29323 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4355
  signal tmp_ivl_29325 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4355
  signal tmp_ivl_2933 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3041
  signal tmp_ivl_29330 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4356
  signal tmp_ivl_29335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4356
  signal tmp_ivl_29337 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4356
  signal tmp_ivl_29342 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4356
  signal tmp_ivl_29344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4356
  signal tmp_ivl_29346 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4356
  signal tmp_ivl_29348 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4356
  signal tmp_ivl_29353 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4357
  signal tmp_ivl_29358 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4357
  signal tmp_ivl_29360 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4357
  signal tmp_ivl_29365 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4357
  signal tmp_ivl_29367 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4357
  signal tmp_ivl_29372 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4358
  signal tmp_ivl_29377 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4358
  signal tmp_ivl_2938 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3041
  signal tmp_ivl_29380 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4358
  signal tmp_ivl_29381 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4358
  signal tmp_ivl_29386 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4358
  signal tmp_ivl_29388 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4358
  signal tmp_ivl_29394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4359
  signal tmp_ivl_29395 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4359
  signal tmp_ivl_294 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2950
  signal tmp_ivl_29400 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4359
  signal tmp_ivl_29403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4359
  signal tmp_ivl_29405 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4359
  signal tmp_ivl_29406 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4359
  signal tmp_ivl_2941 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3041
  signal tmp_ivl_29411 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4359
  signal tmp_ivl_29413 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4359
  signal tmp_ivl_29418 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4360
  signal tmp_ivl_29423 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4360
  signal tmp_ivl_29425 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4360
  signal tmp_ivl_2943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3041
  signal tmp_ivl_29430 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4360
  signal tmp_ivl_29432 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4360
  signal tmp_ivl_29437 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4361
  signal tmp_ivl_2944 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3041
  signal tmp_ivl_29442 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4361
  signal tmp_ivl_29444 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4361
  signal tmp_ivl_29449 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4361
  signal tmp_ivl_29451 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4361
  signal tmp_ivl_29453 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4361
  signal tmp_ivl_29455 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4361
  signal tmp_ivl_29460 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4362
  signal tmp_ivl_29465 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4362
  signal tmp_ivl_29468 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4362
  signal tmp_ivl_29469 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4362
  signal tmp_ivl_29474 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4362
  signal tmp_ivl_29476 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4362
  signal tmp_ivl_29482 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4363
  signal tmp_ivl_29483 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4363
  signal tmp_ivl_29488 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4363
  signal tmp_ivl_2949 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3041
  signal tmp_ivl_29491 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4363
  signal tmp_ivl_29493 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4363
  signal tmp_ivl_29494 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4363
  signal tmp_ivl_29499 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4363
  signal tmp_ivl_29501 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4363
  signal tmp_ivl_29506 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4364
  signal tmp_ivl_2951 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3041
  signal tmp_ivl_29511 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4364
  signal tmp_ivl_29513 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4364
  signal tmp_ivl_29518 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4364
  signal tmp_ivl_29520 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4364
  signal tmp_ivl_29525 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4365
  signal tmp_ivl_2953 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3041
  signal tmp_ivl_29530 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4365
  signal tmp_ivl_29532 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4365
  signal tmp_ivl_29537 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4365
  signal tmp_ivl_29539 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4365
  signal tmp_ivl_29544 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4366
  signal tmp_ivl_29549 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4366
  signal tmp_ivl_29551 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4366
  signal tmp_ivl_29556 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4366
  signal tmp_ivl_29558 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4366
  signal tmp_ivl_29560 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4366
  signal tmp_ivl_29562 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4366
  signal tmp_ivl_29567 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4367
  signal tmp_ivl_29572 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4367
  signal tmp_ivl_29575 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4367
  signal tmp_ivl_29576 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4367
  signal tmp_ivl_29581 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4367
  signal tmp_ivl_29583 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4367
  signal tmp_ivl_29589 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4368
  signal tmp_ivl_2959 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3042
  signal tmp_ivl_29590 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4368
  signal tmp_ivl_29595 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4368
  signal tmp_ivl_29598 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4368
  signal tmp_ivl_29600 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4368
  signal tmp_ivl_29601 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4368
  signal tmp_ivl_29606 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4368
  signal tmp_ivl_29608 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4368
  signal tmp_ivl_2961 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3042
  signal tmp_ivl_29613 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4369
  signal tmp_ivl_29618 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4369
  signal tmp_ivl_2962 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3042
  signal tmp_ivl_29620 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4369
  signal tmp_ivl_29625 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4369
  signal tmp_ivl_29627 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4369
  signal tmp_ivl_29632 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4370
  signal tmp_ivl_29637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4370
  signal tmp_ivl_29639 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4370
  signal tmp_ivl_29644 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4370
  signal tmp_ivl_29646 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4370
  signal tmp_ivl_29651 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4371
  signal tmp_ivl_29656 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4371
  signal tmp_ivl_29658 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4371
  signal tmp_ivl_29663 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4371
  signal tmp_ivl_29665 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4371
  signal tmp_ivl_29667 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4371
  signal tmp_ivl_29669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4371
  signal tmp_ivl_2967 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3042
  signal tmp_ivl_29674 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4372
  signal tmp_ivl_29679 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4372
  signal tmp_ivl_29681 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4372
  signal tmp_ivl_29686 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4372
  signal tmp_ivl_29688 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4372
  signal tmp_ivl_29693 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4373
  signal tmp_ivl_29698 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4373
  signal tmp_ivl_2970 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3042
  signal tmp_ivl_29701 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4373
  signal tmp_ivl_29702 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4373
  signal tmp_ivl_29707 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4373
  signal tmp_ivl_29709 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4373
  signal tmp_ivl_29715 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4374
  signal tmp_ivl_29716 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4374
  signal tmp_ivl_2972 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3042
  signal tmp_ivl_29721 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4374
  signal tmp_ivl_29724 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4374
  signal tmp_ivl_29726 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4374
  signal tmp_ivl_29727 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4374
  signal tmp_ivl_2973 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3042
  signal tmp_ivl_29732 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4374
  signal tmp_ivl_29734 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4374
  signal tmp_ivl_29739 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4375
  signal tmp_ivl_29744 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4375
  signal tmp_ivl_29746 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4375
  signal tmp_ivl_29751 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4375
  signal tmp_ivl_29753 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4375
  signal tmp_ivl_29758 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4376
  signal tmp_ivl_29763 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4376
  signal tmp_ivl_29765 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4376
  signal tmp_ivl_29770 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4376
  signal tmp_ivl_29772 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4376
  signal tmp_ivl_29774 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4376
  signal tmp_ivl_29776 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4376
  signal tmp_ivl_2978 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3042
  signal tmp_ivl_29781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4377
  signal tmp_ivl_29786 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4377
  signal tmp_ivl_29789 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4377
  signal tmp_ivl_29790 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4377
  signal tmp_ivl_29795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4377
  signal tmp_ivl_29797 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4377
  signal tmp_ivl_2980 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3042
  signal tmp_ivl_29803 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4378
  signal tmp_ivl_29804 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4378
  signal tmp_ivl_29809 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4378
  signal tmp_ivl_29812 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4378
  signal tmp_ivl_29814 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4378
  signal tmp_ivl_29815 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4378
  signal tmp_ivl_2982 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3042
  signal tmp_ivl_29820 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4378
  signal tmp_ivl_29822 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4378
  signal tmp_ivl_29827 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4379
  signal tmp_ivl_29832 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4379
  signal tmp_ivl_29834 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4379
  signal tmp_ivl_29839 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4379
  signal tmp_ivl_29841 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4379
  signal tmp_ivl_29846 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4380
  signal tmp_ivl_29851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4380
  signal tmp_ivl_29853 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4380
  signal tmp_ivl_29858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4380
  signal tmp_ivl_29860 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4380
  signal tmp_ivl_29865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4381
  signal tmp_ivl_29870 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4381
  signal tmp_ivl_29872 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4381
  signal tmp_ivl_29877 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4381
  signal tmp_ivl_29879 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4381
  signal tmp_ivl_2988 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3043
  signal tmp_ivl_29881 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4381
  signal tmp_ivl_29883 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4381
  signal tmp_ivl_29888 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4382
  signal tmp_ivl_29893 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4382
  signal tmp_ivl_29896 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4382
  signal tmp_ivl_29897 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4382
  signal tmp_ivl_299 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2950
  signal tmp_ivl_2990 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3043
  signal tmp_ivl_29902 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4382
  signal tmp_ivl_29904 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4382
  signal tmp_ivl_2991 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3043
  signal tmp_ivl_29910 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4383
  signal tmp_ivl_29911 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4383
  signal tmp_ivl_29916 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4383
  signal tmp_ivl_29919 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4383
  signal tmp_ivl_29921 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4383
  signal tmp_ivl_29922 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4383
  signal tmp_ivl_29927 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4383
  signal tmp_ivl_29929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4383
  signal tmp_ivl_29934 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4384
  signal tmp_ivl_29939 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4384
  signal tmp_ivl_29941 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4384
  signal tmp_ivl_29946 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4384
  signal tmp_ivl_29948 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4384
  signal tmp_ivl_29953 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4385
  signal tmp_ivl_29958 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4385
  signal tmp_ivl_2996 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3043
  signal tmp_ivl_29960 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4385
  signal tmp_ivl_29965 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4385
  signal tmp_ivl_29967 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4385
  signal tmp_ivl_29972 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4386
  signal tmp_ivl_29977 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4386
  signal tmp_ivl_29979 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4386
  signal tmp_ivl_29984 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4386
  signal tmp_ivl_29986 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4386
  signal tmp_ivl_29988 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4386
  signal tmp_ivl_2999 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3043
  signal tmp_ivl_29990 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4386
  signal tmp_ivl_29995 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4387
  signal tmp_ivl_3 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2940
  signal tmp_ivl_30 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2941
  signal tmp_ivl_30000 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4387
  signal tmp_ivl_30003 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4387
  signal tmp_ivl_30004 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4387
  signal tmp_ivl_30009 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4387
  signal tmp_ivl_3001 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3043
  signal tmp_ivl_30011 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4387
  signal tmp_ivl_30017 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4388
  signal tmp_ivl_30018 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4388
  signal tmp_ivl_3002 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3043
  signal tmp_ivl_30023 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4388
  signal tmp_ivl_30026 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4388
  signal tmp_ivl_30028 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4388
  signal tmp_ivl_30029 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4388
  signal tmp_ivl_30034 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4388
  signal tmp_ivl_30036 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4388
  signal tmp_ivl_30041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4389
  signal tmp_ivl_30046 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4389
  signal tmp_ivl_30048 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4389
  signal tmp_ivl_30053 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4389
  signal tmp_ivl_30055 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4389
  signal tmp_ivl_30060 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4390
  signal tmp_ivl_30065 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4390
  signal tmp_ivl_30067 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4390
  signal tmp_ivl_3007 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3043
  signal tmp_ivl_30072 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4390
  signal tmp_ivl_30074 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4390
  signal tmp_ivl_30079 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4391
  signal tmp_ivl_30084 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4391
  signal tmp_ivl_30086 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4391
  signal tmp_ivl_3009 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3043
  signal tmp_ivl_30091 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4391
  signal tmp_ivl_30093 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4391
  signal tmp_ivl_30095 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4391
  signal tmp_ivl_30097 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4391
  signal tmp_ivl_30102 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4392
  signal tmp_ivl_30107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4392
  signal tmp_ivl_3011 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3043
  signal tmp_ivl_30110 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4392
  signal tmp_ivl_30111 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4392
  signal tmp_ivl_30116 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4392
  signal tmp_ivl_30118 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4392
  signal tmp_ivl_30124 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4393
  signal tmp_ivl_30125 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4393
  signal tmp_ivl_30130 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4393
  signal tmp_ivl_30133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4393
  signal tmp_ivl_30135 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4393
  signal tmp_ivl_30136 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4393
  signal tmp_ivl_30141 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4393
  signal tmp_ivl_30143 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4393
  signal tmp_ivl_30148 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4394
  signal tmp_ivl_30153 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4394
  signal tmp_ivl_30155 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4394
  signal tmp_ivl_30160 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4394
  signal tmp_ivl_30162 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4394
  signal tmp_ivl_30167 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4395
  signal tmp_ivl_3017 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3044
  signal tmp_ivl_30172 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4395
  signal tmp_ivl_30174 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4395
  signal tmp_ivl_30179 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4395
  signal tmp_ivl_30181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4395
  signal tmp_ivl_30186 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4396
  signal tmp_ivl_3019 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3044
  signal tmp_ivl_30191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4396
  signal tmp_ivl_30193 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4396
  signal tmp_ivl_30198 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4396
  signal tmp_ivl_302 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2950
  signal tmp_ivl_3020 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3044
  signal tmp_ivl_30200 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4396
  signal tmp_ivl_30202 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4396
  signal tmp_ivl_30204 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4396
  signal tmp_ivl_30209 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4397
  signal tmp_ivl_30214 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4397
  signal tmp_ivl_30217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4397
  signal tmp_ivl_30218 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4397
  signal tmp_ivl_30223 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4397
  signal tmp_ivl_30225 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4397
  signal tmp_ivl_30231 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4398
  signal tmp_ivl_30232 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4398
  signal tmp_ivl_30237 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4398
  signal tmp_ivl_30240 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4398
  signal tmp_ivl_30242 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4398
  signal tmp_ivl_30243 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4398
  signal tmp_ivl_30248 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4398
  signal tmp_ivl_3025 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3044
  signal tmp_ivl_30250 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4398
  signal tmp_ivl_30255 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4399
  signal tmp_ivl_30260 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4399
  signal tmp_ivl_30262 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4399
  signal tmp_ivl_30267 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4399
  signal tmp_ivl_30269 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4399
  signal tmp_ivl_30274 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4400
  signal tmp_ivl_30279 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4400
  signal tmp_ivl_3028 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3044
  signal tmp_ivl_30281 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4400
  signal tmp_ivl_30286 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4400
  signal tmp_ivl_30288 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4400
  signal tmp_ivl_30293 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4401
  signal tmp_ivl_30298 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4401
  signal tmp_ivl_3030 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3044
  signal tmp_ivl_30300 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4401
  signal tmp_ivl_30305 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4401
  signal tmp_ivl_30307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4401
  signal tmp_ivl_30309 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4401
  signal tmp_ivl_3031 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3044
  signal tmp_ivl_30311 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4401
  signal tmp_ivl_30317 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4402
  signal tmp_ivl_30318 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4402
  signal tmp_ivl_30323 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4402
  signal tmp_ivl_30325 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4402
  signal tmp_ivl_30330 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4402
  signal tmp_ivl_30332 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4402
  signal tmp_ivl_30337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4403
  signal tmp_ivl_30340 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4403
  signal tmp_ivl_30341 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4403
  signal tmp_ivl_30346 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4403
  signal tmp_ivl_30348 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4403
  signal tmp_ivl_30353 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4403
  signal tmp_ivl_30355 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4403
  signal tmp_ivl_3036 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3044
  signal tmp_ivl_30360 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4404
  signal tmp_ivl_30365 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4404
  signal tmp_ivl_30368 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4404
  signal tmp_ivl_30369 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4404
  signal tmp_ivl_30374 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4404
  signal tmp_ivl_30376 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4404
  signal tmp_ivl_3038 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3044
  signal tmp_ivl_30381 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4405
  signal tmp_ivl_30386 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4405
  signal tmp_ivl_30389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4405
  signal tmp_ivl_30391 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4405
  signal tmp_ivl_30392 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4405
  signal tmp_ivl_30397 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4405
  signal tmp_ivl_30399 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4405
  signal tmp_ivl_304 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2950
  signal tmp_ivl_3040 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3044
  signal tmp_ivl_30404 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4406
  signal tmp_ivl_30409 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4406
  signal tmp_ivl_30411 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4406
  signal tmp_ivl_30416 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4406
  signal tmp_ivl_30418 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4406
  signal tmp_ivl_30423 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4407
  signal tmp_ivl_30428 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4407
  signal tmp_ivl_30430 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4407
  signal tmp_ivl_30435 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4407
  signal tmp_ivl_30437 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4407
  signal tmp_ivl_30439 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4407
  signal tmp_ivl_30441 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4407
  signal tmp_ivl_30446 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4408
  signal tmp_ivl_30451 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4408
  signal tmp_ivl_30453 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4408
  signal tmp_ivl_30458 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4408
  signal tmp_ivl_3046 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3045
  signal tmp_ivl_30460 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4408
  signal tmp_ivl_30465 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4409
  signal tmp_ivl_30470 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4409
  signal tmp_ivl_30472 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4409
  signal tmp_ivl_30477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4409
  signal tmp_ivl_30479 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4409
  signal tmp_ivl_3048 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3045
  signal tmp_ivl_30481 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4409
  signal tmp_ivl_30483 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4409
  signal tmp_ivl_30488 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4410
  signal tmp_ivl_3049 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3045
  signal tmp_ivl_30493 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4410
  signal tmp_ivl_30496 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4410
  signal tmp_ivl_30497 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4410
  signal tmp_ivl_305 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2950
  signal tmp_ivl_30502 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4410
  signal tmp_ivl_30504 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4410
  signal tmp_ivl_30510 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4411
  signal tmp_ivl_30511 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4411
  signal tmp_ivl_30516 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4411
  signal tmp_ivl_30519 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4411
  signal tmp_ivl_30521 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4411
  signal tmp_ivl_30522 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4411
  signal tmp_ivl_30527 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4411
  signal tmp_ivl_30529 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4411
  signal tmp_ivl_30534 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4412
  signal tmp_ivl_30539 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4412
  signal tmp_ivl_3054 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3045
  signal tmp_ivl_30541 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4412
  signal tmp_ivl_30546 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4412
  signal tmp_ivl_30548 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4412
  signal tmp_ivl_30553 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4413
  signal tmp_ivl_30558 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4413
  signal tmp_ivl_30560 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4413
  signal tmp_ivl_30565 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4413
  signal tmp_ivl_30567 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4413
  signal tmp_ivl_3057 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3045
  signal tmp_ivl_30572 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4414
  signal tmp_ivl_30577 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4414
  signal tmp_ivl_30579 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4414
  signal tmp_ivl_30584 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4414
  signal tmp_ivl_30586 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4414
  signal tmp_ivl_30588 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4414
  signal tmp_ivl_3059 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3045
  signal tmp_ivl_30590 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4414
  signal tmp_ivl_30595 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4415
  signal tmp_ivl_3060 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3045
  signal tmp_ivl_30600 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4415
  signal tmp_ivl_30603 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4415
  signal tmp_ivl_30604 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4415
  signal tmp_ivl_30609 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4415
  signal tmp_ivl_30611 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4415
  signal tmp_ivl_30617 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4416
  signal tmp_ivl_30618 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4416
  signal tmp_ivl_30623 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4416
  signal tmp_ivl_30626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4416
  signal tmp_ivl_30628 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4416
  signal tmp_ivl_30629 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4416
  signal tmp_ivl_30634 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4416
  signal tmp_ivl_30636 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4416
  signal tmp_ivl_30641 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4417
  signal tmp_ivl_30646 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4417
  signal tmp_ivl_30648 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4417
  signal tmp_ivl_3065 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3045
  signal tmp_ivl_30653 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4417
  signal tmp_ivl_30655 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4417
  signal tmp_ivl_30660 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4418
  signal tmp_ivl_30665 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4418
  signal tmp_ivl_30667 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4418
  signal tmp_ivl_3067 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3045
  signal tmp_ivl_30672 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4418
  signal tmp_ivl_30674 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4418
  signal tmp_ivl_30679 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4419
  signal tmp_ivl_30684 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4419
  signal tmp_ivl_30686 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4419
  signal tmp_ivl_3069 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3045
  signal tmp_ivl_30691 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4419
  signal tmp_ivl_30693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4419
  signal tmp_ivl_30695 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4419
  signal tmp_ivl_30697 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4419
  signal tmp_ivl_30702 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4420
  signal tmp_ivl_30707 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4420
  signal tmp_ivl_30710 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4420
  signal tmp_ivl_30711 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4420
  signal tmp_ivl_30716 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4420
  signal tmp_ivl_30718 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4420
  signal tmp_ivl_30723 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4421
  signal tmp_ivl_30728 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4421
  signal tmp_ivl_30731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4421
  signal tmp_ivl_30732 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4421
  signal tmp_ivl_30737 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4421
  signal tmp_ivl_30739 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4421
  signal tmp_ivl_30744 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4422
  signal tmp_ivl_30749 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4422
  signal tmp_ivl_3075 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3046
  signal tmp_ivl_30752 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4422
  signal tmp_ivl_30754 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4422
  signal tmp_ivl_30755 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4422
  signal tmp_ivl_30760 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4422
  signal tmp_ivl_30762 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4422
  signal tmp_ivl_30767 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4423
  signal tmp_ivl_3077 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3046
  signal tmp_ivl_30772 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4423
  signal tmp_ivl_30774 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4423
  signal tmp_ivl_30779 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4423
  signal tmp_ivl_3078 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3046
  signal tmp_ivl_30781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4423
  signal tmp_ivl_30786 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4424
  signal tmp_ivl_30791 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4424
  signal tmp_ivl_30793 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4424
  signal tmp_ivl_30798 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4424
  signal tmp_ivl_30800 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4424
  signal tmp_ivl_30802 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4424
  signal tmp_ivl_30804 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4424
  signal tmp_ivl_30809 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4425
  signal tmp_ivl_30814 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4425
  signal tmp_ivl_30816 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4425
  signal tmp_ivl_30821 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4425
  signal tmp_ivl_30823 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4425
  signal tmp_ivl_30828 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4426
  signal tmp_ivl_3083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3046
  signal tmp_ivl_30833 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4426
  signal tmp_ivl_30835 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4426
  signal tmp_ivl_30840 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4426
  signal tmp_ivl_30842 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4426
  signal tmp_ivl_30844 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4426
  signal tmp_ivl_30846 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4426
  signal tmp_ivl_30852 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4427
  signal tmp_ivl_30853 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4427
  signal tmp_ivl_30858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4427
  signal tmp_ivl_3086 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3046
  signal tmp_ivl_30860 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4427
  signal tmp_ivl_30865 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4427
  signal tmp_ivl_30867 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4427
  signal tmp_ivl_30872 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4428
  signal tmp_ivl_30877 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4428
  signal tmp_ivl_3088 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3046
  signal tmp_ivl_30880 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4428
  signal tmp_ivl_30881 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4428
  signal tmp_ivl_30886 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4428
  signal tmp_ivl_30888 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4428
  signal tmp_ivl_3089 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3046
  signal tmp_ivl_30893 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4429
  signal tmp_ivl_30898 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4429
  signal tmp_ivl_30900 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4429
  signal tmp_ivl_30905 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4429
  signal tmp_ivl_30907 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4429
  signal tmp_ivl_30912 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4430
  signal tmp_ivl_30917 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4430
  signal tmp_ivl_30919 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4430
  signal tmp_ivl_30924 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4430
  signal tmp_ivl_30926 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4430
  signal tmp_ivl_30928 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4430
  signal tmp_ivl_30930 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4430
  signal tmp_ivl_30935 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4431
  signal tmp_ivl_3094 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3046
  signal tmp_ivl_30940 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4431
  signal tmp_ivl_30942 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4431
  signal tmp_ivl_30947 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4431
  signal tmp_ivl_30949 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4431
  signal tmp_ivl_30955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4432
  signal tmp_ivl_30956 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4432
  signal tmp_ivl_3096 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3046
  signal tmp_ivl_30961 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4432
  signal tmp_ivl_30964 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4432
  signal tmp_ivl_30966 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4432
  signal tmp_ivl_30967 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4432
  signal tmp_ivl_30972 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4432
  signal tmp_ivl_30974 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4432
  signal tmp_ivl_30979 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4433
  signal tmp_ivl_3098 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3046
  signal tmp_ivl_30984 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4433
  signal tmp_ivl_30986 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4433
  signal tmp_ivl_30991 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4433
  signal tmp_ivl_30993 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4433
  signal tmp_ivl_30998 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4434
  signal tmp_ivl_310 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2950
  signal tmp_ivl_31003 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4434
  signal tmp_ivl_31005 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4434
  signal tmp_ivl_31010 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4434
  signal tmp_ivl_31012 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4434
  signal tmp_ivl_31014 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4434
  signal tmp_ivl_31016 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4434
  signal tmp_ivl_31021 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4435
  signal tmp_ivl_31026 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4435
  signal tmp_ivl_31028 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4435
  signal tmp_ivl_31033 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4435
  signal tmp_ivl_31035 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4435
  signal tmp_ivl_3104 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3047
  signal tmp_ivl_31040 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4436
  signal tmp_ivl_31045 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4436
  signal tmp_ivl_31047 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4436
  signal tmp_ivl_31052 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4436
  signal tmp_ivl_31054 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4436
  signal tmp_ivl_31056 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4436
  signal tmp_ivl_31058 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4436
  signal tmp_ivl_3106 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3047
  signal tmp_ivl_31064 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4437
  signal tmp_ivl_31065 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4437
  signal tmp_ivl_3107 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3047
  signal tmp_ivl_31070 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4437
  signal tmp_ivl_31072 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4437
  signal tmp_ivl_31077 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4437
  signal tmp_ivl_31079 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4437
  signal tmp_ivl_31084 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4438
  signal tmp_ivl_31086 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4438
  signal tmp_ivl_31091 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4438
  signal tmp_ivl_31093 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4438
  signal tmp_ivl_31098 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4438
  signal tmp_ivl_31100 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4438
  signal tmp_ivl_31105 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4439
  signal tmp_ivl_31110 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4439
  signal tmp_ivl_31113 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4439
  signal tmp_ivl_31114 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4439
  signal tmp_ivl_31119 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4439
  signal tmp_ivl_3112 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3047
  signal tmp_ivl_31121 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4439
  signal tmp_ivl_31127 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4440
  signal tmp_ivl_31129 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4440
  signal tmp_ivl_31130 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4440
  signal tmp_ivl_31135 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4440
  signal tmp_ivl_31137 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4440
  signal tmp_ivl_31142 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4440
  signal tmp_ivl_31144 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4440
  signal tmp_ivl_31149 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4441
  signal tmp_ivl_3115 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3047
  signal tmp_ivl_31154 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4441
  signal tmp_ivl_31156 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4441
  signal tmp_ivl_31161 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4441
  signal tmp_ivl_31163 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4441
  signal tmp_ivl_31168 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4442
  signal tmp_ivl_3117 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3047
  signal tmp_ivl_31173 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4442
  signal tmp_ivl_31175 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4442
  signal tmp_ivl_3118 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3047
  signal tmp_ivl_31180 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4442
  signal tmp_ivl_31182 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4442
  signal tmp_ivl_31184 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4442
  signal tmp_ivl_31186 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4442
  signal tmp_ivl_31191 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4443
  signal tmp_ivl_31196 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4443
  signal tmp_ivl_31198 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4443
  signal tmp_ivl_312 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2950
  signal tmp_ivl_31203 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4443
  signal tmp_ivl_31205 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4443
  signal tmp_ivl_31210 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4444
  signal tmp_ivl_31215 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4444
  signal tmp_ivl_31217 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4444
  signal tmp_ivl_31222 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4444
  signal tmp_ivl_31224 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4444
  signal tmp_ivl_31226 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4444
  signal tmp_ivl_31228 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4444
  signal tmp_ivl_3123 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3047
  signal tmp_ivl_31233 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4445
  signal tmp_ivl_31238 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4445
  signal tmp_ivl_31240 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4445
  signal tmp_ivl_31245 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4445
  signal tmp_ivl_31247 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4445
  signal tmp_ivl_3125 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3047
  signal tmp_ivl_31252 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4446
  signal tmp_ivl_31257 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4446
  signal tmp_ivl_31259 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4446
  signal tmp_ivl_31264 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4446
  signal tmp_ivl_31266 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4446
  signal tmp_ivl_31268 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4446
  signal tmp_ivl_3127 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3047
  signal tmp_ivl_31270 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4446
  signal tmp_ivl_31276 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4447
  signal tmp_ivl_31277 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4447
  signal tmp_ivl_31282 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4447
  signal tmp_ivl_31284 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4447
  signal tmp_ivl_31289 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4447
  signal tmp_ivl_31291 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4447
  signal tmp_ivl_31297 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4448
  signal tmp_ivl_31298 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4448
  signal tmp_ivl_31303 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4448
  signal tmp_ivl_31306 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4448
  signal tmp_ivl_31308 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4448
  signal tmp_ivl_31309 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4448
  signal tmp_ivl_31314 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4448
  signal tmp_ivl_31316 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4448
  signal tmp_ivl_31321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4449
  signal tmp_ivl_31326 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4449
  signal tmp_ivl_31328 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4449
  signal tmp_ivl_3133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3048
  signal tmp_ivl_31333 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4449
  signal tmp_ivl_31335 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4449
  signal tmp_ivl_31340 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4450
  signal tmp_ivl_31345 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4450
  signal tmp_ivl_31347 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4450
  signal tmp_ivl_3135 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3048
  signal tmp_ivl_31352 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4450
  signal tmp_ivl_31354 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4450
  signal tmp_ivl_31359 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4451
  signal tmp_ivl_3136 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3048
  signal tmp_ivl_31364 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4451
  signal tmp_ivl_31366 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4451
  signal tmp_ivl_31371 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4451
  signal tmp_ivl_31373 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4451
  signal tmp_ivl_31375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4451
  signal tmp_ivl_31377 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4451
  signal tmp_ivl_31382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4452
  signal tmp_ivl_31387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4452
  signal tmp_ivl_31389 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4452
  signal tmp_ivl_31394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4452
  signal tmp_ivl_31396 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4452
  signal tmp_ivl_314 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2950
  signal tmp_ivl_31401 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4453
  signal tmp_ivl_31406 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4453
  signal tmp_ivl_31408 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4453
  signal tmp_ivl_3141 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3048
  signal tmp_ivl_31413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4453
  signal tmp_ivl_31415 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4453
  signal tmp_ivl_31417 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4453
  signal tmp_ivl_31419 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4453
  signal tmp_ivl_31424 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4454
  signal tmp_ivl_31429 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4454
  signal tmp_ivl_31431 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4454
  signal tmp_ivl_31436 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4454
  signal tmp_ivl_31438 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4454
  signal tmp_ivl_3144 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3048
  signal tmp_ivl_31443 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4455
  signal tmp_ivl_31448 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4455
  signal tmp_ivl_31450 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4455
  signal tmp_ivl_31455 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4455
  signal tmp_ivl_31457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4455
  signal tmp_ivl_31459 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4455
  signal tmp_ivl_3146 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3048
  signal tmp_ivl_31461 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4455
  signal tmp_ivl_31467 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4456
  signal tmp_ivl_31468 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4456
  signal tmp_ivl_3147 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3048
  signal tmp_ivl_31473 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4456
  signal tmp_ivl_31475 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4456
  signal tmp_ivl_31480 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4456
  signal tmp_ivl_31482 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4456
  signal tmp_ivl_31487 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4457
  signal tmp_ivl_31492 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4457
  signal tmp_ivl_31494 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4457
  signal tmp_ivl_31499 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4457
  signal tmp_ivl_31501 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4457
  signal tmp_ivl_31506 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4458
  signal tmp_ivl_31511 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4458
  signal tmp_ivl_31513 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4458
  signal tmp_ivl_31518 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4458
  signal tmp_ivl_3152 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3048
  signal tmp_ivl_31520 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4458
  signal tmp_ivl_31522 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4458
  signal tmp_ivl_31524 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4458
  signal tmp_ivl_31529 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4459
  signal tmp_ivl_31534 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4459
  signal tmp_ivl_31536 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4459
  signal tmp_ivl_3154 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3048
  signal tmp_ivl_31541 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4459
  signal tmp_ivl_31543 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4459
  signal tmp_ivl_31548 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4460
  signal tmp_ivl_31553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4460
  signal tmp_ivl_31555 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4460
  signal tmp_ivl_3156 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3048
  signal tmp_ivl_31560 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4460
  signal tmp_ivl_31562 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4460
  signal tmp_ivl_31564 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4460
  signal tmp_ivl_31566 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4460
  signal tmp_ivl_31571 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4461
  signal tmp_ivl_31576 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4461
  signal tmp_ivl_31579 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4461
  signal tmp_ivl_31580 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4461
  signal tmp_ivl_31585 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4461
  signal tmp_ivl_31587 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4461
  signal tmp_ivl_31592 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4462
  signal tmp_ivl_31597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4462
  signal tmp_ivl_31599 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4462
  signal tmp_ivl_31604 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4462
  signal tmp_ivl_31606 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4462
  signal tmp_ivl_31611 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4463
  signal tmp_ivl_31616 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4463
  signal tmp_ivl_31619 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4463
  signal tmp_ivl_3162 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3049
  signal tmp_ivl_31620 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4463
  signal tmp_ivl_31625 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4463
  signal tmp_ivl_31627 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4463
  signal tmp_ivl_31632 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4464
  signal tmp_ivl_31637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4464
  signal tmp_ivl_31639 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4464
  signal tmp_ivl_3164 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3049
  signal tmp_ivl_31644 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4464
  signal tmp_ivl_31646 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4464
  signal tmp_ivl_31648 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4464
  signal tmp_ivl_3165 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3049
  signal tmp_ivl_31650 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4464
  signal tmp_ivl_31656 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4465
  signal tmp_ivl_31657 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4465
  signal tmp_ivl_31662 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4465
  signal tmp_ivl_31665 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4465
  signal tmp_ivl_31667 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4465
  signal tmp_ivl_31668 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4465
  signal tmp_ivl_31673 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4465
  signal tmp_ivl_31675 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4465
  signal tmp_ivl_31680 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4466
  signal tmp_ivl_31685 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4466
  signal tmp_ivl_31687 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4466
  signal tmp_ivl_31692 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4466
  signal tmp_ivl_31694 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4466
  signal tmp_ivl_31699 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4467
  signal tmp_ivl_3170 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3049
  signal tmp_ivl_31704 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4467
  signal tmp_ivl_31706 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4467
  signal tmp_ivl_31711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4467
  signal tmp_ivl_31713 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4467
  signal tmp_ivl_31718 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4468
  signal tmp_ivl_31723 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4468
  signal tmp_ivl_31725 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4468
  signal tmp_ivl_3173 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3049
  signal tmp_ivl_31730 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4468
  signal tmp_ivl_31732 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4468
  signal tmp_ivl_31734 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4468
  signal tmp_ivl_31736 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4468
  signal tmp_ivl_31741 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4469
  signal tmp_ivl_31746 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4469
  signal tmp_ivl_31748 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4469
  signal tmp_ivl_3175 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3049
  signal tmp_ivl_31753 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4469
  signal tmp_ivl_31755 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4469
  signal tmp_ivl_3176 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3049
  signal tmp_ivl_31760 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4470
  signal tmp_ivl_31765 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4470
  signal tmp_ivl_31767 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4470
  signal tmp_ivl_31772 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4470
  signal tmp_ivl_31774 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4470
  signal tmp_ivl_31776 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4470
  signal tmp_ivl_31778 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4470
  signal tmp_ivl_31783 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4471
  signal tmp_ivl_31788 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4471
  signal tmp_ivl_31790 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4471
  signal tmp_ivl_31795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4471
  signal tmp_ivl_31797 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4471
  signal tmp_ivl_31802 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4472
  signal tmp_ivl_31807 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4472
  signal tmp_ivl_31809 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4472
  signal tmp_ivl_3181 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3049
  signal tmp_ivl_31814 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4472
  signal tmp_ivl_31816 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4472
  signal tmp_ivl_31818 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4472
  signal tmp_ivl_31820 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4472
  signal tmp_ivl_31825 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4473
  signal tmp_ivl_3183 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3049
  signal tmp_ivl_31830 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4473
  signal tmp_ivl_31832 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4473
  signal tmp_ivl_31837 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4473
  signal tmp_ivl_31839 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4473
  signal tmp_ivl_31845 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4474
  signal tmp_ivl_31846 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4474
  signal tmp_ivl_3185 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3049
  signal tmp_ivl_31851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4474
  signal tmp_ivl_31853 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4474
  signal tmp_ivl_31858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4474
  signal tmp_ivl_31860 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4474
  signal tmp_ivl_31865 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4475
  signal tmp_ivl_31868 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4475
  signal tmp_ivl_31869 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4475
  signal tmp_ivl_31874 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4475
  signal tmp_ivl_31876 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4475
  signal tmp_ivl_31881 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4475
  signal tmp_ivl_31883 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4475
  signal tmp_ivl_31888 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4476
  signal tmp_ivl_31893 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4476
  signal tmp_ivl_31895 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4476
  signal tmp_ivl_31900 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4476
  signal tmp_ivl_31902 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4476
  signal tmp_ivl_31904 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4476
  signal tmp_ivl_31906 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4476
  signal tmp_ivl_3191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3050
  signal tmp_ivl_31911 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4477
  signal tmp_ivl_31916 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4477
  signal tmp_ivl_31918 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4477
  signal tmp_ivl_31923 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4477
  signal tmp_ivl_31925 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4477
  signal tmp_ivl_3193 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3050
  signal tmp_ivl_31930 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4478
  signal tmp_ivl_31935 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4478
  signal tmp_ivl_31937 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4478
  signal tmp_ivl_3194 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3050
  signal tmp_ivl_31942 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4478
  signal tmp_ivl_31944 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4478
  signal tmp_ivl_31949 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4479
  signal tmp_ivl_31952 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4479
  signal tmp_ivl_31953 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4479
  signal tmp_ivl_31958 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4479
  signal tmp_ivl_31960 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4479
  signal tmp_ivl_31965 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4479
  signal tmp_ivl_31967 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4479
  signal tmp_ivl_31969 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4479
  signal tmp_ivl_31971 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4479
  signal tmp_ivl_31976 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4480
  signal tmp_ivl_31981 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4480
  signal tmp_ivl_31983 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4480
  signal tmp_ivl_31988 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4480
  signal tmp_ivl_3199 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3050
  signal tmp_ivl_31990 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4480
  signal tmp_ivl_31995 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4481
  signal tmp_ivl_32 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2941
  signal tmp_ivl_320 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2951
  signal tmp_ivl_32000 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4481
  signal tmp_ivl_32002 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4481
  signal tmp_ivl_32007 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4481
  signal tmp_ivl_32009 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4481
  signal tmp_ivl_32011 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4481
  signal tmp_ivl_32013 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4481
  signal tmp_ivl_32018 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4482
  signal tmp_ivl_3202 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3050
  signal tmp_ivl_32023 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4482
  signal tmp_ivl_32025 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4482
  signal tmp_ivl_32030 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4482
  signal tmp_ivl_32032 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4482
  signal tmp_ivl_32037 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4483
  signal tmp_ivl_3204 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3050
  signal tmp_ivl_32042 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4483
  signal tmp_ivl_32044 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4483
  signal tmp_ivl_32049 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4483
  signal tmp_ivl_3205 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3050
  signal tmp_ivl_32051 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4483
  signal tmp_ivl_32053 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4483
  signal tmp_ivl_32055 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4483
  signal tmp_ivl_32060 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4484
  signal tmp_ivl_32065 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4484
  signal tmp_ivl_32067 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4484
  signal tmp_ivl_32072 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4484
  signal tmp_ivl_32074 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4484
  signal tmp_ivl_32079 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4485
  signal tmp_ivl_32084 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4485
  signal tmp_ivl_32086 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4485
  signal tmp_ivl_32091 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4485
  signal tmp_ivl_32093 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4485
  signal tmp_ivl_32095 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4485
  signal tmp_ivl_32097 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4485
  signal tmp_ivl_3210 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3050
  signal tmp_ivl_32102 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4486
  signal tmp_ivl_32107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4486
  signal tmp_ivl_32109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4486
  signal tmp_ivl_32114 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4486
  signal tmp_ivl_32116 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4486
  signal tmp_ivl_3212 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3050
  signal tmp_ivl_32121 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4487
  signal tmp_ivl_32126 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4487
  signal tmp_ivl_32128 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4487
  signal tmp_ivl_32133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4487
  signal tmp_ivl_32135 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4487
  signal tmp_ivl_32137 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4487
  signal tmp_ivl_32139 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4487
  signal tmp_ivl_3214 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3050
  signal tmp_ivl_32144 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4488
  signal tmp_ivl_32149 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4488
  signal tmp_ivl_32151 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4488
  signal tmp_ivl_32156 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4488
  signal tmp_ivl_32158 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4488
  signal tmp_ivl_32163 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4489
  signal tmp_ivl_32168 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4489
  signal tmp_ivl_32170 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4489
  signal tmp_ivl_32175 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4489
  signal tmp_ivl_32177 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4489
  signal tmp_ivl_32179 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4489
  signal tmp_ivl_32181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4489
  signal tmp_ivl_32186 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4490
  signal tmp_ivl_32191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4490
  signal tmp_ivl_32193 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4490
  signal tmp_ivl_32198 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4490
  signal tmp_ivl_322 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2951
  signal tmp_ivl_3220 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3051
  signal tmp_ivl_32200 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4490
  signal tmp_ivl_32205 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4491
  signal tmp_ivl_32210 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4491
  signal tmp_ivl_32212 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4491
  signal tmp_ivl_32217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4491
  signal tmp_ivl_32219 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4491
  signal tmp_ivl_3222 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3051
  signal tmp_ivl_32221 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4491
  signal tmp_ivl_32223 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4491
  signal tmp_ivl_32228 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4492
  signal tmp_ivl_3223 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3051
  signal tmp_ivl_32233 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4492
  signal tmp_ivl_32235 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4492
  signal tmp_ivl_32240 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4492
  signal tmp_ivl_32242 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4492
  signal tmp_ivl_32247 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4493
  signal tmp_ivl_32252 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4493
  signal tmp_ivl_32254 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4493
  signal tmp_ivl_32259 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4493
  signal tmp_ivl_32261 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4493
  signal tmp_ivl_32263 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4493
  signal tmp_ivl_32265 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4493
  signal tmp_ivl_32270 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4494
  signal tmp_ivl_32275 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4494
  signal tmp_ivl_32277 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4494
  signal tmp_ivl_3228 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3051
  signal tmp_ivl_32282 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4494
  signal tmp_ivl_32284 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4494
  signal tmp_ivl_32289 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4495
  signal tmp_ivl_32294 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4495
  signal tmp_ivl_32296 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4495
  signal tmp_ivl_323 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2951
  signal tmp_ivl_32301 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4495
  signal tmp_ivl_32303 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4495
  signal tmp_ivl_32305 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4495
  signal tmp_ivl_32307 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4495
  signal tmp_ivl_3231 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3051
  signal tmp_ivl_32312 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4496
  signal tmp_ivl_32317 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4496
  signal tmp_ivl_32319 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4496
  signal tmp_ivl_32324 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4496
  signal tmp_ivl_32326 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4496
  signal tmp_ivl_3233 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3051
  signal tmp_ivl_32331 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4497
  signal tmp_ivl_32336 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4497
  signal tmp_ivl_32338 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4497
  signal tmp_ivl_3234 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3051
  signal tmp_ivl_32343 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4497
  signal tmp_ivl_32345 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4497
  signal tmp_ivl_32347 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4497
  signal tmp_ivl_32349 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4497
  signal tmp_ivl_32354 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4498
  signal tmp_ivl_32359 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4498
  signal tmp_ivl_32361 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4498
  signal tmp_ivl_32366 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4498
  signal tmp_ivl_32368 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4498
  signal tmp_ivl_32373 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4499
  signal tmp_ivl_32378 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4499
  signal tmp_ivl_32380 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4499
  signal tmp_ivl_32385 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4499
  signal tmp_ivl_32387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4499
  signal tmp_ivl_32389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4499
  signal tmp_ivl_3239 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3051
  signal tmp_ivl_32391 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4499
  signal tmp_ivl_32396 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4500
  signal tmp_ivl_32401 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4500
  signal tmp_ivl_32403 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4500
  signal tmp_ivl_32408 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4500
  signal tmp_ivl_3241 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3051
  signal tmp_ivl_32410 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4500
  signal tmp_ivl_32415 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4501
  signal tmp_ivl_32420 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4501
  signal tmp_ivl_32422 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4501
  signal tmp_ivl_32427 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4501
  signal tmp_ivl_32429 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4501
  signal tmp_ivl_3243 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3051
  signal tmp_ivl_32431 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4501
  signal tmp_ivl_32433 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4501
  signal tmp_ivl_32438 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4502
  signal tmp_ivl_32443 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4502
  signal tmp_ivl_32445 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4502
  signal tmp_ivl_32450 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4502
  signal tmp_ivl_32452 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4502
  signal tmp_ivl_32457 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4503
  signal tmp_ivl_32462 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4503
  signal tmp_ivl_32464 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4503
  signal tmp_ivl_32469 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4503
  signal tmp_ivl_32471 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4503
  signal tmp_ivl_32473 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4503
  signal tmp_ivl_32475 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4503
  signal tmp_ivl_32480 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4504
  signal tmp_ivl_32485 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4504
  signal tmp_ivl_32487 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4504
  signal tmp_ivl_3249 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3052
  signal tmp_ivl_32492 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4504
  signal tmp_ivl_32494 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4504
  signal tmp_ivl_32499 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4505
  signal tmp_ivl_32504 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4505
  signal tmp_ivl_32506 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4505
  signal tmp_ivl_3251 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3052
  signal tmp_ivl_32511 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4505
  signal tmp_ivl_32513 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4505
  signal tmp_ivl_32515 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4505
  signal tmp_ivl_32517 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4505
  signal tmp_ivl_3252 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3052
  signal tmp_ivl_32522 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4506
  signal tmp_ivl_32527 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4506
  signal tmp_ivl_32529 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4506
  signal tmp_ivl_32534 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4506
  signal tmp_ivl_32536 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4506
  signal tmp_ivl_32541 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4507
  signal tmp_ivl_32546 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4507
  signal tmp_ivl_32548 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4507
  signal tmp_ivl_32553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4507
  signal tmp_ivl_32555 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4507
  signal tmp_ivl_32557 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4507
  signal tmp_ivl_32559 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4507
  signal tmp_ivl_32564 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4508
  signal tmp_ivl_32569 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4508
  signal tmp_ivl_3257 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3052
  signal tmp_ivl_32571 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4508
  signal tmp_ivl_32576 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4508
  signal tmp_ivl_32578 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4508
  signal tmp_ivl_32583 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4509
  signal tmp_ivl_32588 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4509
  signal tmp_ivl_32590 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4509
  signal tmp_ivl_32595 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4509
  signal tmp_ivl_32597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4509
  signal tmp_ivl_32599 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4509
  signal tmp_ivl_3260 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3052
  signal tmp_ivl_32601 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4509
  signal tmp_ivl_32606 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4510
  signal tmp_ivl_32611 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4510
  signal tmp_ivl_32613 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4510
  signal tmp_ivl_32618 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4510
  signal tmp_ivl_3262 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3052
  signal tmp_ivl_32620 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4510
  signal tmp_ivl_32625 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4511
  signal tmp_ivl_3263 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3052
  signal tmp_ivl_32630 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4511
  signal tmp_ivl_32632 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4511
  signal tmp_ivl_32637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4511
  signal tmp_ivl_32639 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4511
  signal tmp_ivl_32641 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4511
  signal tmp_ivl_32643 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4511
  signal tmp_ivl_32648 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4512
  signal tmp_ivl_32653 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4512
  signal tmp_ivl_32655 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4512
  signal tmp_ivl_32660 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4512
  signal tmp_ivl_32662 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4512
  signal tmp_ivl_32667 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4513
  signal tmp_ivl_32672 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4513
  signal tmp_ivl_32674 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4513
  signal tmp_ivl_32679 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4513
  signal tmp_ivl_3268 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3052
  signal tmp_ivl_32681 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4513
  signal tmp_ivl_32683 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4513
  signal tmp_ivl_32685 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4513
  signal tmp_ivl_32690 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4514
  signal tmp_ivl_32695 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4514
  signal tmp_ivl_32697 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4514
  signal tmp_ivl_3270 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3052
  signal tmp_ivl_32702 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4514
  signal tmp_ivl_32704 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4514
  signal tmp_ivl_32709 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4515
  signal tmp_ivl_32714 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4515
  signal tmp_ivl_32716 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4515
  signal tmp_ivl_3272 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3052
  signal tmp_ivl_32721 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4515
  signal tmp_ivl_32723 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4515
  signal tmp_ivl_32725 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4515
  signal tmp_ivl_32727 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4515
  signal tmp_ivl_32732 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4516
  signal tmp_ivl_32737 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4516
  signal tmp_ivl_32739 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4516
  signal tmp_ivl_32744 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4516
  signal tmp_ivl_32746 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4516
  signal tmp_ivl_32751 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4517
  signal tmp_ivl_32756 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4517
  signal tmp_ivl_32758 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4517
  signal tmp_ivl_32763 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4517
  signal tmp_ivl_32765 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4517
  signal tmp_ivl_32767 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4517
  signal tmp_ivl_32769 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4517
  signal tmp_ivl_32774 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4518
  signal tmp_ivl_32779 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4518
  signal tmp_ivl_3278 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3053
  signal tmp_ivl_32781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4518
  signal tmp_ivl_32786 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4518
  signal tmp_ivl_32788 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4518
  signal tmp_ivl_32793 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4519
  signal tmp_ivl_32798 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4519
  signal tmp_ivl_328 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2951
  signal tmp_ivl_3280 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3053
  signal tmp_ivl_32800 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4519
  signal tmp_ivl_32805 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4519
  signal tmp_ivl_32807 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4519
  signal tmp_ivl_32809 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4519
  signal tmp_ivl_3281 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3053
  signal tmp_ivl_32811 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4519
  signal tmp_ivl_32816 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4520
  signal tmp_ivl_32821 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4520
  signal tmp_ivl_32823 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4520
  signal tmp_ivl_32828 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4520
  signal tmp_ivl_32830 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4520
  signal tmp_ivl_32835 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4521
  signal tmp_ivl_32840 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4521
  signal tmp_ivl_32842 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4521
  signal tmp_ivl_32847 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4521
  signal tmp_ivl_32849 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4521
  signal tmp_ivl_32851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4521
  signal tmp_ivl_32853 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4521
  signal tmp_ivl_32858 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4522
  signal tmp_ivl_3286 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3053
  signal tmp_ivl_32863 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4522
  signal tmp_ivl_32865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4522
  signal tmp_ivl_32870 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4522
  signal tmp_ivl_32872 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4522
  signal tmp_ivl_32877 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4523
  signal tmp_ivl_32882 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4523
  signal tmp_ivl_32884 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4523
  signal tmp_ivl_32889 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4523
  signal tmp_ivl_3289 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3053
  signal tmp_ivl_32891 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4523
  signal tmp_ivl_32893 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4523
  signal tmp_ivl_32895 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4523
  signal tmp_ivl_32900 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4524
  signal tmp_ivl_32905 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4524
  signal tmp_ivl_32907 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4524
  signal tmp_ivl_3291 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3053
  signal tmp_ivl_32912 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4524
  signal tmp_ivl_32914 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4524
  signal tmp_ivl_32919 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4525
  signal tmp_ivl_3292 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3053
  signal tmp_ivl_32924 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4525
  signal tmp_ivl_32926 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4525
  signal tmp_ivl_32931 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4525
  signal tmp_ivl_32933 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4525
  signal tmp_ivl_32935 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4525
  signal tmp_ivl_32937 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4525
  signal tmp_ivl_32942 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4526
  signal tmp_ivl_32947 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4526
  signal tmp_ivl_32949 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4526
  signal tmp_ivl_32954 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4526
  signal tmp_ivl_32956 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4526
  signal tmp_ivl_32961 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4527
  signal tmp_ivl_32966 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4527
  signal tmp_ivl_32968 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4527
  signal tmp_ivl_3297 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3053
  signal tmp_ivl_32973 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4527
  signal tmp_ivl_32975 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4527
  signal tmp_ivl_32977 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4527
  signal tmp_ivl_32979 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4527
  signal tmp_ivl_32984 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4528
  signal tmp_ivl_32989 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4528
  signal tmp_ivl_3299 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3053
  signal tmp_ivl_32991 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4528
  signal tmp_ivl_32996 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4528
  signal tmp_ivl_32998 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4528
  signal tmp_ivl_33 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2941
  signal tmp_ivl_33003 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4529
  signal tmp_ivl_33008 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4529
  signal tmp_ivl_3301 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3053
  signal tmp_ivl_33010 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4529
  signal tmp_ivl_33015 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4529
  signal tmp_ivl_33017 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4529
  signal tmp_ivl_33019 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4529
  signal tmp_ivl_33021 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4529
  signal tmp_ivl_33026 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4530
  signal tmp_ivl_33031 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4530
  signal tmp_ivl_33033 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4530
  signal tmp_ivl_33038 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4530
  signal tmp_ivl_33040 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4530
  signal tmp_ivl_33045 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4531
  signal tmp_ivl_33050 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4531
  signal tmp_ivl_33052 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4531
  signal tmp_ivl_33057 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4531
  signal tmp_ivl_33059 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4531
  signal tmp_ivl_33061 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4531
  signal tmp_ivl_33063 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4531
  signal tmp_ivl_33068 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4532
  signal tmp_ivl_3307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3054
  signal tmp_ivl_33073 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4532
  signal tmp_ivl_33075 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4532
  signal tmp_ivl_33080 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4532
  signal tmp_ivl_33082 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4532
  signal tmp_ivl_33087 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4533
  signal tmp_ivl_3309 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3054
  signal tmp_ivl_33092 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4533
  signal tmp_ivl_33094 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4533
  signal tmp_ivl_33099 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4533
  signal tmp_ivl_331 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2951
  signal tmp_ivl_3310 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3054
  signal tmp_ivl_33101 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4533
  signal tmp_ivl_33103 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4533
  signal tmp_ivl_33105 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4533
  signal tmp_ivl_33110 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4534
  signal tmp_ivl_33115 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4534
  signal tmp_ivl_33117 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4534
  signal tmp_ivl_33122 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4534
  signal tmp_ivl_33124 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4534
  signal tmp_ivl_33129 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4535
  signal tmp_ivl_33134 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4535
  signal tmp_ivl_33136 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4535
  signal tmp_ivl_33141 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4535
  signal tmp_ivl_33143 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4535
  signal tmp_ivl_33145 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4535
  signal tmp_ivl_33147 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4535
  signal tmp_ivl_3315 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3054
  signal tmp_ivl_33152 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4536
  signal tmp_ivl_33157 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4536
  signal tmp_ivl_33159 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4536
  signal tmp_ivl_33164 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4536
  signal tmp_ivl_33166 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4536
  signal tmp_ivl_33171 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4537
  signal tmp_ivl_33176 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4537
  signal tmp_ivl_33178 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4537
  signal tmp_ivl_3318 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3054
  signal tmp_ivl_33183 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4537
  signal tmp_ivl_33185 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4537
  signal tmp_ivl_33187 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4537
  signal tmp_ivl_33189 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4537
  signal tmp_ivl_33194 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4538
  signal tmp_ivl_33199 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4538
  signal tmp_ivl_3320 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3054
  signal tmp_ivl_33201 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4538
  signal tmp_ivl_33206 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4538
  signal tmp_ivl_33208 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4538
  signal tmp_ivl_3321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3054
  signal tmp_ivl_33213 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4539
  signal tmp_ivl_33218 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4539
  signal tmp_ivl_33220 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4539
  signal tmp_ivl_33225 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4539
  signal tmp_ivl_33227 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4539
  signal tmp_ivl_33229 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4539
  signal tmp_ivl_33231 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4539
  signal tmp_ivl_33236 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4540
  signal tmp_ivl_33241 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4540
  signal tmp_ivl_33243 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4540
  signal tmp_ivl_33248 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4540
  signal tmp_ivl_33250 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4540
  signal tmp_ivl_33255 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4541
  signal tmp_ivl_3326 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3054
  signal tmp_ivl_33260 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4541
  signal tmp_ivl_33262 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4541
  signal tmp_ivl_33267 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4541
  signal tmp_ivl_33269 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4541
  signal tmp_ivl_33271 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4541
  signal tmp_ivl_33273 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4541
  signal tmp_ivl_33278 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4542
  signal tmp_ivl_3328 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3054
  signal tmp_ivl_33283 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4542
  signal tmp_ivl_33285 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4542
  signal tmp_ivl_33290 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4542
  signal tmp_ivl_33292 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4542
  signal tmp_ivl_33297 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4543
  signal tmp_ivl_333 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2951
  signal tmp_ivl_3330 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3054
  signal tmp_ivl_33302 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4543
  signal tmp_ivl_33304 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4543
  signal tmp_ivl_33309 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4543
  signal tmp_ivl_33311 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4543
  signal tmp_ivl_33313 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4543
  signal tmp_ivl_33315 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4543
  signal tmp_ivl_33320 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4544
  signal tmp_ivl_33325 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4544
  signal tmp_ivl_33327 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4544
  signal tmp_ivl_33332 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4544
  signal tmp_ivl_33334 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4544
  signal tmp_ivl_33339 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4545
  signal tmp_ivl_33344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4545
  signal tmp_ivl_33346 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4545
  signal tmp_ivl_33351 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4545
  signal tmp_ivl_33353 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4545
  signal tmp_ivl_33355 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4545
  signal tmp_ivl_33357 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4545
  signal tmp_ivl_3336 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3055
  signal tmp_ivl_33362 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4546
  signal tmp_ivl_33367 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4546
  signal tmp_ivl_33369 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4546
  signal tmp_ivl_33374 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4546
  signal tmp_ivl_33376 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4546
  signal tmp_ivl_3338 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3055
  signal tmp_ivl_33381 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4547
  signal tmp_ivl_33386 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4547
  signal tmp_ivl_33388 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4547
  signal tmp_ivl_3339 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3055
  signal tmp_ivl_33393 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4547
  signal tmp_ivl_33395 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4547
  signal tmp_ivl_33397 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4547
  signal tmp_ivl_33399 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4547
  signal tmp_ivl_334 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2951
  signal tmp_ivl_33404 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4548
  signal tmp_ivl_33409 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4548
  signal tmp_ivl_33411 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4548
  signal tmp_ivl_33416 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4548
  signal tmp_ivl_33418 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4548
  signal tmp_ivl_33423 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4549
  signal tmp_ivl_33428 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4549
  signal tmp_ivl_33430 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4549
  signal tmp_ivl_33435 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4549
  signal tmp_ivl_33437 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4549
  signal tmp_ivl_33439 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4549
  signal tmp_ivl_3344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3055
  signal tmp_ivl_33441 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4549
  signal tmp_ivl_33446 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4550
  signal tmp_ivl_33451 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4550
  signal tmp_ivl_33453 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4550
  signal tmp_ivl_33458 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4550
  signal tmp_ivl_33460 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4550
  signal tmp_ivl_33465 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4551
  signal tmp_ivl_3347 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3055
  signal tmp_ivl_33470 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4551
  signal tmp_ivl_33472 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4551
  signal tmp_ivl_33477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4551
  signal tmp_ivl_33479 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4551
  signal tmp_ivl_33481 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4551
  signal tmp_ivl_33483 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4551
  signal tmp_ivl_33488 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4552
  signal tmp_ivl_3349 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3055
  signal tmp_ivl_33493 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4552
  signal tmp_ivl_33495 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4552
  signal tmp_ivl_3350 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3055
  signal tmp_ivl_33500 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4552
  signal tmp_ivl_33502 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4552
  signal tmp_ivl_33507 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4553
  signal tmp_ivl_33512 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4553
  signal tmp_ivl_33514 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4553
  signal tmp_ivl_33519 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4553
  signal tmp_ivl_33521 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4553
  signal tmp_ivl_33523 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4553
  signal tmp_ivl_33525 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4553
  signal tmp_ivl_33530 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4554
  signal tmp_ivl_33535 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4554
  signal tmp_ivl_33537 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4554
  signal tmp_ivl_33542 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4554
  signal tmp_ivl_33544 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4554
  signal tmp_ivl_33549 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4555
  signal tmp_ivl_3355 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3055
  signal tmp_ivl_33554 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4555
  signal tmp_ivl_33556 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4555
  signal tmp_ivl_33561 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4555
  signal tmp_ivl_33563 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4555
  signal tmp_ivl_33565 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4555
  signal tmp_ivl_33567 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4555
  signal tmp_ivl_3357 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3055
  signal tmp_ivl_33572 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4556
  signal tmp_ivl_33577 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4556
  signal tmp_ivl_33579 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4556
  signal tmp_ivl_33584 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4556
  signal tmp_ivl_33586 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4556
  signal tmp_ivl_3359 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3055
  signal tmp_ivl_33591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4557
  signal tmp_ivl_33596 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4557
  signal tmp_ivl_33598 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4557
  signal tmp_ivl_33603 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4557
  signal tmp_ivl_33605 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4557
  signal tmp_ivl_33607 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4557
  signal tmp_ivl_33609 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4557
  signal tmp_ivl_33614 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4558
  signal tmp_ivl_33619 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4558
  signal tmp_ivl_33621 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4558
  signal tmp_ivl_33626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4558
  signal tmp_ivl_33628 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4558
  signal tmp_ivl_33633 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4559
  signal tmp_ivl_33638 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4559
  signal tmp_ivl_33640 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4559
  signal tmp_ivl_33645 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4559
  signal tmp_ivl_33647 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4559
  signal tmp_ivl_33649 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4559
  signal tmp_ivl_3365 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3056
  signal tmp_ivl_33651 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4559
  signal tmp_ivl_33656 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4560
  signal tmp_ivl_33661 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4560
  signal tmp_ivl_33663 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4560
  signal tmp_ivl_33668 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4560
  signal tmp_ivl_3367 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3056
  signal tmp_ivl_33670 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4560
  signal tmp_ivl_33675 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4561
  signal tmp_ivl_3368 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3056
  signal tmp_ivl_33680 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4561
  signal tmp_ivl_33682 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4561
  signal tmp_ivl_33687 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4561
  signal tmp_ivl_33689 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4561
  signal tmp_ivl_33691 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4561
  signal tmp_ivl_33693 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4561
  signal tmp_ivl_33698 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4562
  signal tmp_ivl_33703 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4562
  signal tmp_ivl_33705 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4562
  signal tmp_ivl_33710 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4562
  signal tmp_ivl_33712 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4562
  signal tmp_ivl_33717 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4563
  signal tmp_ivl_33722 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4563
  signal tmp_ivl_33724 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4563
  signal tmp_ivl_33729 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4563
  signal tmp_ivl_3373 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3056
  signal tmp_ivl_33731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4563
  signal tmp_ivl_33733 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4563
  signal tmp_ivl_33735 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4563
  signal tmp_ivl_33740 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4564
  signal tmp_ivl_33745 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4564
  signal tmp_ivl_33747 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4564
  signal tmp_ivl_33752 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4564
  signal tmp_ivl_33754 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4564
  signal tmp_ivl_33759 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4565
  signal tmp_ivl_3376 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3056
  signal tmp_ivl_33764 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4565
  signal tmp_ivl_33766 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4565
  signal tmp_ivl_33771 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4565
  signal tmp_ivl_33773 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4565
  signal tmp_ivl_33775 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4565
  signal tmp_ivl_33777 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4565
  signal tmp_ivl_3378 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3056
  signal tmp_ivl_33782 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4566
  signal tmp_ivl_33787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4566
  signal tmp_ivl_33789 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4566
  signal tmp_ivl_3379 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3056
  signal tmp_ivl_33794 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4566
  signal tmp_ivl_33796 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4566
  signal tmp_ivl_33801 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4567
  signal tmp_ivl_33806 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4567
  signal tmp_ivl_33808 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4567
  signal tmp_ivl_33813 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4567
  signal tmp_ivl_33815 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4567
  signal tmp_ivl_33817 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4567
  signal tmp_ivl_33819 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4567
  signal tmp_ivl_33824 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4568
  signal tmp_ivl_33829 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4568
  signal tmp_ivl_33831 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4568
  signal tmp_ivl_33836 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4568
  signal tmp_ivl_33838 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4568
  signal tmp_ivl_3384 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3056
  signal tmp_ivl_33843 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4569
  signal tmp_ivl_33848 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4569
  signal tmp_ivl_33850 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4569
  signal tmp_ivl_33855 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4569
  signal tmp_ivl_33857 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4569
  signal tmp_ivl_33859 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4569
  signal tmp_ivl_3386 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3056
  signal tmp_ivl_33861 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4569
  signal tmp_ivl_33866 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4570
  signal tmp_ivl_33871 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4570
  signal tmp_ivl_33873 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4570
  signal tmp_ivl_33878 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4570
  signal tmp_ivl_3388 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3056
  signal tmp_ivl_33880 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4570
  signal tmp_ivl_33885 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4571
  signal tmp_ivl_33890 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4571
  signal tmp_ivl_33892 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4571
  signal tmp_ivl_33897 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4571
  signal tmp_ivl_33899 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4571
  signal tmp_ivl_339 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2951
  signal tmp_ivl_33901 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4571
  signal tmp_ivl_33903 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4571
  signal tmp_ivl_33908 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4572
  signal tmp_ivl_33913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4572
  signal tmp_ivl_33915 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4572
  signal tmp_ivl_33920 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4572
  signal tmp_ivl_33922 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4572
  signal tmp_ivl_33927 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4573
  signal tmp_ivl_33932 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4573
  signal tmp_ivl_33934 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4573
  signal tmp_ivl_33939 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4573
  signal tmp_ivl_3394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3057
  signal tmp_ivl_33941 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4573
  signal tmp_ivl_33943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4573
  signal tmp_ivl_33945 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4573
  signal tmp_ivl_33950 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4574
  signal tmp_ivl_33955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4574
  signal tmp_ivl_33957 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4574
  signal tmp_ivl_3396 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3057
  signal tmp_ivl_33962 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4574
  signal tmp_ivl_33964 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4574
  signal tmp_ivl_33969 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4575
  signal tmp_ivl_3397 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3057
  signal tmp_ivl_33974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4575
  signal tmp_ivl_33976 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4575
  signal tmp_ivl_33981 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4575
  signal tmp_ivl_33983 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4575
  signal tmp_ivl_33985 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4575
  signal tmp_ivl_33987 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4575
  signal tmp_ivl_33992 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4576
  signal tmp_ivl_33997 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4576
  signal tmp_ivl_33999 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4576
  signal tmp_ivl_34004 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4576
  signal tmp_ivl_34006 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4576
  signal tmp_ivl_34011 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4577
  signal tmp_ivl_34016 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4577
  signal tmp_ivl_34018 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4577
  signal tmp_ivl_3402 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3057
  signal tmp_ivl_34023 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4577
  signal tmp_ivl_34025 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4577
  signal tmp_ivl_34027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4577
  signal tmp_ivl_34029 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4577
  signal tmp_ivl_34034 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4578
  signal tmp_ivl_34039 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4578
  signal tmp_ivl_34041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4578
  signal tmp_ivl_34046 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4578
  signal tmp_ivl_34048 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4578
  signal tmp_ivl_3405 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3057
  signal tmp_ivl_34053 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4579
  signal tmp_ivl_34058 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4579
  signal tmp_ivl_34060 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4579
  signal tmp_ivl_34065 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4579
  signal tmp_ivl_34067 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4579
  signal tmp_ivl_34069 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4579
  signal tmp_ivl_3407 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3057
  signal tmp_ivl_34071 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4579
  signal tmp_ivl_34076 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4580
  signal tmp_ivl_3408 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3057
  signal tmp_ivl_34081 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4580
  signal tmp_ivl_34083 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4580
  signal tmp_ivl_34088 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4580
  signal tmp_ivl_34090 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4580
  signal tmp_ivl_34095 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4581
  signal tmp_ivl_341 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2951
  signal tmp_ivl_34100 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4581
  signal tmp_ivl_34102 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4581
  signal tmp_ivl_34107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4581
  signal tmp_ivl_34109 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4581
  signal tmp_ivl_34111 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4581
  signal tmp_ivl_34113 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4581
  signal tmp_ivl_34118 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4582
  signal tmp_ivl_34123 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4582
  signal tmp_ivl_34125 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4582
  signal tmp_ivl_3413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3057
  signal tmp_ivl_34130 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4582
  signal tmp_ivl_34132 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4582
  signal tmp_ivl_34137 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4583
  signal tmp_ivl_34139 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4583
  signal tmp_ivl_34144 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4583
  signal tmp_ivl_34146 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4583
  signal tmp_ivl_3415 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3057
  signal tmp_ivl_34151 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4583
  signal tmp_ivl_34153 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4583
  signal tmp_ivl_34158 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4584
  signal tmp_ivl_34163 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4584
  signal tmp_ivl_34165 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4584
  signal tmp_ivl_3417 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3057
  signal tmp_ivl_34170 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4584
  signal tmp_ivl_34172 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4584
  signal tmp_ivl_34174 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4584
  signal tmp_ivl_34176 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4584
  signal tmp_ivl_34181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4585
  signal tmp_ivl_34186 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4585
  signal tmp_ivl_34189 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4585
  signal tmp_ivl_34190 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4585
  signal tmp_ivl_34195 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4585
  signal tmp_ivl_34197 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4585
  signal tmp_ivl_34202 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4586
  signal tmp_ivl_34207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4586
  signal tmp_ivl_34209 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4586
  signal tmp_ivl_34214 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4586
  signal tmp_ivl_34216 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4586
  signal tmp_ivl_34221 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4587
  signal tmp_ivl_34226 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4587
  signal tmp_ivl_34228 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4587
  signal tmp_ivl_3423 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3058
  signal tmp_ivl_34233 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4587
  signal tmp_ivl_34235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4587
  signal tmp_ivl_34237 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4587
  signal tmp_ivl_34239 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4587
  signal tmp_ivl_34244 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4588
  signal tmp_ivl_34249 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4588
  signal tmp_ivl_3425 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3058
  signal tmp_ivl_34251 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4588
  signal tmp_ivl_34256 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4588
  signal tmp_ivl_34258 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4588
  signal tmp_ivl_3426 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3058
  signal tmp_ivl_34263 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4589
  signal tmp_ivl_34268 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4589
  signal tmp_ivl_34270 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4589
  signal tmp_ivl_34275 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4589
  signal tmp_ivl_34277 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4589
  signal tmp_ivl_34279 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4589
  signal tmp_ivl_34281 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4589
  signal tmp_ivl_34286 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4590
  signal tmp_ivl_34291 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4590
  signal tmp_ivl_34293 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4590
  signal tmp_ivl_34298 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4590
  signal tmp_ivl_343 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2951
  signal tmp_ivl_34300 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4590
  signal tmp_ivl_34305 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4591
  signal tmp_ivl_3431 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3058
  signal tmp_ivl_34310 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4591
  signal tmp_ivl_34312 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4591
  signal tmp_ivl_34317 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4591
  signal tmp_ivl_34319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4591
  signal tmp_ivl_34321 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4591
  signal tmp_ivl_34323 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4591
  signal tmp_ivl_34328 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4592
  signal tmp_ivl_34333 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4592
  signal tmp_ivl_34335 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4592
  signal tmp_ivl_3434 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3058
  signal tmp_ivl_34340 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4592
  signal tmp_ivl_34342 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4592
  signal tmp_ivl_34347 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4593
  signal tmp_ivl_34352 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4593
  signal tmp_ivl_34354 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4593
  signal tmp_ivl_34359 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4593
  signal tmp_ivl_3436 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3058
  signal tmp_ivl_34361 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4593
  signal tmp_ivl_34363 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4593
  signal tmp_ivl_34365 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4593
  signal tmp_ivl_3437 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3058
  signal tmp_ivl_34370 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4594
  signal tmp_ivl_34375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4594
  signal tmp_ivl_34377 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4594
  signal tmp_ivl_34382 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4594
  signal tmp_ivl_34384 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4594
  signal tmp_ivl_34389 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4595
  signal tmp_ivl_34394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4595
  signal tmp_ivl_34396 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4595
  signal tmp_ivl_34401 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4595
  signal tmp_ivl_34403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4595
  signal tmp_ivl_34405 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4595
  signal tmp_ivl_34407 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4595
  signal tmp_ivl_34412 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4596
  signal tmp_ivl_34417 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4596
  signal tmp_ivl_34419 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4596
  signal tmp_ivl_3442 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3058
  signal tmp_ivl_34424 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4596
  signal tmp_ivl_34426 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4596
  signal tmp_ivl_34431 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4597
  signal tmp_ivl_34436 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4597
  signal tmp_ivl_34438 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4597
  signal tmp_ivl_3444 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3058
  signal tmp_ivl_34443 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4597
  signal tmp_ivl_34445 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4597
  signal tmp_ivl_34447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4597
  signal tmp_ivl_34449 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4597
  signal tmp_ivl_34455 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4598
  signal tmp_ivl_34456 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4598
  signal tmp_ivl_3446 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3058
  signal tmp_ivl_34461 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4598
  signal tmp_ivl_34464 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4598
  signal tmp_ivl_34466 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4598
  signal tmp_ivl_34467 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4598
  signal tmp_ivl_34472 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4598
  signal tmp_ivl_34474 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4598
  signal tmp_ivl_34479 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4599
  signal tmp_ivl_34484 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4599
  signal tmp_ivl_34486 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4599
  signal tmp_ivl_34491 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4599
  signal tmp_ivl_34493 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4599
  signal tmp_ivl_34498 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4600
  signal tmp_ivl_34503 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4600
  signal tmp_ivl_34505 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4600
  signal tmp_ivl_34510 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4600
  signal tmp_ivl_34512 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4600
  signal tmp_ivl_34517 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4601
  signal tmp_ivl_3452 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3059
  signal tmp_ivl_34522 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4601
  signal tmp_ivl_34524 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4601
  signal tmp_ivl_34529 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4601
  signal tmp_ivl_34531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4601
  signal tmp_ivl_34533 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4601
  signal tmp_ivl_34535 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4601
  signal tmp_ivl_3454 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3059
  signal tmp_ivl_34540 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4602
  signal tmp_ivl_34545 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4602
  signal tmp_ivl_34547 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4602
  signal tmp_ivl_3455 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3059
  signal tmp_ivl_34552 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4602
  signal tmp_ivl_34554 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4602
  signal tmp_ivl_34559 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4603
  signal tmp_ivl_34564 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4603
  signal tmp_ivl_34566 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4603
  signal tmp_ivl_34571 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4603
  signal tmp_ivl_34573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4603
  signal tmp_ivl_34575 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4603
  signal tmp_ivl_34577 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4603
  signal tmp_ivl_34582 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4604
  signal tmp_ivl_34587 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4604
  signal tmp_ivl_34589 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4604
  signal tmp_ivl_34594 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4604
  signal tmp_ivl_34596 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4604
  signal tmp_ivl_3460 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3059
  signal tmp_ivl_34601 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4605
  signal tmp_ivl_34606 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4605
  signal tmp_ivl_34608 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4605
  signal tmp_ivl_34613 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4605
  signal tmp_ivl_34615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4605
  signal tmp_ivl_34617 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4605
  signal tmp_ivl_34619 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4605
  signal tmp_ivl_34625 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4606
  signal tmp_ivl_34626 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4606
  signal tmp_ivl_3463 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3059
  signal tmp_ivl_34631 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4606
  signal tmp_ivl_34634 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4606
  signal tmp_ivl_34636 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4606
  signal tmp_ivl_34637 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4606
  signal tmp_ivl_34642 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4606
  signal tmp_ivl_34644 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4606
  signal tmp_ivl_34649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4607
  signal tmp_ivl_3465 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3059
  signal tmp_ivl_34654 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4607
  signal tmp_ivl_34656 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4607
  signal tmp_ivl_3466 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3059
  signal tmp_ivl_34661 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4607
  signal tmp_ivl_34663 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4607
  signal tmp_ivl_34668 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4608
  signal tmp_ivl_34673 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4608
  signal tmp_ivl_34675 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4608
  signal tmp_ivl_34680 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4608
  signal tmp_ivl_34682 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4608
  signal tmp_ivl_34687 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4609
  signal tmp_ivl_34692 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4609
  signal tmp_ivl_34694 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4609
  signal tmp_ivl_34699 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4609
  signal tmp_ivl_34701 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4609
  signal tmp_ivl_34703 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4609
  signal tmp_ivl_34705 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4609
  signal tmp_ivl_3471 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3059
  signal tmp_ivl_34710 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4610
  signal tmp_ivl_34715 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4610
  signal tmp_ivl_34717 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4610
  signal tmp_ivl_34722 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4610
  signal tmp_ivl_34724 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4610
  signal tmp_ivl_34729 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4611
  signal tmp_ivl_3473 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3059
  signal tmp_ivl_34734 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4611
  signal tmp_ivl_34736 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4611
  signal tmp_ivl_34741 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4611
  signal tmp_ivl_34743 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4611
  signal tmp_ivl_34745 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4611
  signal tmp_ivl_34747 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4611
  signal tmp_ivl_3475 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3059
  signal tmp_ivl_34752 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4612
  signal tmp_ivl_34757 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4612
  signal tmp_ivl_34759 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4612
  signal tmp_ivl_34764 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4612
  signal tmp_ivl_34766 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4612
  signal tmp_ivl_34771 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4613
  signal tmp_ivl_34776 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4613
  signal tmp_ivl_34778 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4613
  signal tmp_ivl_34783 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4613
  signal tmp_ivl_34785 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4613
  signal tmp_ivl_34787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4613
  signal tmp_ivl_34789 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4613
  signal tmp_ivl_34795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4614
  signal tmp_ivl_34796 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4614
  signal tmp_ivl_34801 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4614
  signal tmp_ivl_34804 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4614
  signal tmp_ivl_34806 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4614
  signal tmp_ivl_34807 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4614
  signal tmp_ivl_3481 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3060
  signal tmp_ivl_34812 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4614
  signal tmp_ivl_34814 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4614
  signal tmp_ivl_34819 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4615
  signal tmp_ivl_34824 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4615
  signal tmp_ivl_34826 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4615
  signal tmp_ivl_3483 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3060
  signal tmp_ivl_34831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4615
  signal tmp_ivl_34833 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4615
  signal tmp_ivl_34838 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4616
  signal tmp_ivl_3484 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3060
  signal tmp_ivl_34843 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4616
  signal tmp_ivl_34845 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4616
  signal tmp_ivl_34850 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4616
  signal tmp_ivl_34852 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4616
  signal tmp_ivl_34857 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4617
  signal tmp_ivl_34862 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4617
  signal tmp_ivl_34864 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4617
  signal tmp_ivl_34869 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4617
  signal tmp_ivl_34871 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4617
  signal tmp_ivl_34873 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4617
  signal tmp_ivl_34875 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4617
  signal tmp_ivl_34880 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4618
  signal tmp_ivl_34885 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4618
  signal tmp_ivl_34887 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4618
  signal tmp_ivl_3489 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3060
  signal tmp_ivl_34892 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4618
  signal tmp_ivl_34894 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4618
  signal tmp_ivl_34899 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4619
  signal tmp_ivl_349 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2952
  signal tmp_ivl_34904 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4619
  signal tmp_ivl_34906 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4619
  signal tmp_ivl_34911 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4619
  signal tmp_ivl_34913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4619
  signal tmp_ivl_34915 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4619
  signal tmp_ivl_34917 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4619
  signal tmp_ivl_3492 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3060
  signal tmp_ivl_34922 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4620
  signal tmp_ivl_34927 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4620
  signal tmp_ivl_34929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4620
  signal tmp_ivl_34934 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4620
  signal tmp_ivl_34936 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4620
  signal tmp_ivl_3494 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3060
  signal tmp_ivl_34941 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4621
  signal tmp_ivl_34946 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4621
  signal tmp_ivl_34948 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4621
  signal tmp_ivl_3495 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3060
  signal tmp_ivl_34953 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4621
  signal tmp_ivl_34955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4621
  signal tmp_ivl_34957 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4621
  signal tmp_ivl_34959 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4621
  signal tmp_ivl_34965 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4622
  signal tmp_ivl_34966 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4622
  signal tmp_ivl_34971 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4622
  signal tmp_ivl_34974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4622
  signal tmp_ivl_34976 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4622
  signal tmp_ivl_34977 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4622
  signal tmp_ivl_34982 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4622
  signal tmp_ivl_34984 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4622
  signal tmp_ivl_34989 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4623
  signal tmp_ivl_34994 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4623
  signal tmp_ivl_34996 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4623
  signal tmp_ivl_3500 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3060
  signal tmp_ivl_35001 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4623
  signal tmp_ivl_35003 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4623
  signal tmp_ivl_35008 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4624
  signal tmp_ivl_35013 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4624
  signal tmp_ivl_35015 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4624
  signal tmp_ivl_3502 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3060
  signal tmp_ivl_35020 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4624
  signal tmp_ivl_35022 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4624
  signal tmp_ivl_35027 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4625
  signal tmp_ivl_35032 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4625
  signal tmp_ivl_35034 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4625
  signal tmp_ivl_35039 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4625
  signal tmp_ivl_3504 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3060
  signal tmp_ivl_35041 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4625
  signal tmp_ivl_35043 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4625
  signal tmp_ivl_35045 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4625
  signal tmp_ivl_35050 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4626
  signal tmp_ivl_35055 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4626
  signal tmp_ivl_35057 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4626
  signal tmp_ivl_35062 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4626
  signal tmp_ivl_35064 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4626
  signal tmp_ivl_35069 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4627
  signal tmp_ivl_35074 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4627
  signal tmp_ivl_35076 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4627
  signal tmp_ivl_35081 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4627
  signal tmp_ivl_35083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4627
  signal tmp_ivl_35085 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4627
  signal tmp_ivl_35087 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4627
  signal tmp_ivl_35092 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4628
  signal tmp_ivl_35097 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4628
  signal tmp_ivl_35099 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4628
  signal tmp_ivl_351 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2952
  signal tmp_ivl_3510 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3061
  signal tmp_ivl_35104 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4628
  signal tmp_ivl_35106 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4628
  signal tmp_ivl_35111 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4629
  signal tmp_ivl_35116 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4629
  signal tmp_ivl_35118 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4629
  signal tmp_ivl_3512 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3061
  signal tmp_ivl_35123 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4629
  signal tmp_ivl_35125 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4629
  signal tmp_ivl_35127 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4629
  signal tmp_ivl_35129 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4629
  signal tmp_ivl_3513 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3061
  signal tmp_ivl_35135 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4630
  signal tmp_ivl_35136 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4630
  signal tmp_ivl_35141 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4630
  signal tmp_ivl_35143 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4630
  signal tmp_ivl_35148 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4630
  signal tmp_ivl_35151 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4630
  signal tmp_ivl_35155 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4630
  signal tmp_ivl_35157 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4630
  signal tmp_ivl_35159 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4630
  signal tmp_ivl_35164 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4631
  signal tmp_ivl_35169 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4631
  signal tmp_ivl_35171 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4631
  signal tmp_ivl_35176 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4631
  signal tmp_ivl_35179 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4631
  signal tmp_ivl_3518 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3061
  signal tmp_ivl_35183 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4631
  signal tmp_ivl_35185 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4631
  signal tmp_ivl_35187 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4631
  signal tmp_ivl_35192 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4632
  signal tmp_ivl_35197 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4632
  signal tmp_ivl_35199 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4632
  signal tmp_ivl_352 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2952
  signal tmp_ivl_35204 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4632
  signal tmp_ivl_35207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4632
  signal tmp_ivl_3521 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3061
  signal tmp_ivl_35211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4632
  signal tmp_ivl_35213 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4632
  signal tmp_ivl_35215 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4632
  signal tmp_ivl_35220 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4633
  signal tmp_ivl_35225 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4633
  signal tmp_ivl_35227 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4633
  signal tmp_ivl_3523 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3061
  signal tmp_ivl_35232 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4633
  signal tmp_ivl_35235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4633
  signal tmp_ivl_35239 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4633
  signal tmp_ivl_3524 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3061
  signal tmp_ivl_35241 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4633
  signal tmp_ivl_35243 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4633
  signal tmp_ivl_35248 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4634
  signal tmp_ivl_35253 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4634
  signal tmp_ivl_35255 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4634
  signal tmp_ivl_35260 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4634
  signal tmp_ivl_35263 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4634
  signal tmp_ivl_35267 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4634
  signal tmp_ivl_35269 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4634
  signal tmp_ivl_35271 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4634
  signal tmp_ivl_35276 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4635
  signal tmp_ivl_35281 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4635
  signal tmp_ivl_35283 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4635
  signal tmp_ivl_35288 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4635
  signal tmp_ivl_3529 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3061
  signal tmp_ivl_35291 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4635
  signal tmp_ivl_35295 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4635
  signal tmp_ivl_35297 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4635
  signal tmp_ivl_35299 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4635
  signal tmp_ivl_35304 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4636
  signal tmp_ivl_35309 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4636
  signal tmp_ivl_3531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3061
  signal tmp_ivl_35311 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4636
  signal tmp_ivl_35316 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4636
  signal tmp_ivl_35319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4636
  signal tmp_ivl_35323 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4636
  signal tmp_ivl_35325 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4636
  signal tmp_ivl_35327 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4636
  signal tmp_ivl_3533 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3061
  signal tmp_ivl_35332 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4637
  signal tmp_ivl_35337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4637
  signal tmp_ivl_35339 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4637
  signal tmp_ivl_35344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4637
  signal tmp_ivl_35347 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4637
  signal tmp_ivl_35351 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4637
  signal tmp_ivl_35353 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4637
  signal tmp_ivl_35355 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4637
  signal tmp_ivl_35360 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4638
  signal tmp_ivl_35365 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4638
  signal tmp_ivl_35367 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4638
  signal tmp_ivl_35372 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4638
  signal tmp_ivl_35375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4638
  signal tmp_ivl_35379 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4638
  signal tmp_ivl_35381 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4638
  signal tmp_ivl_35383 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4638
  signal tmp_ivl_35388 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4639
  signal tmp_ivl_3539 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3062
  signal tmp_ivl_35393 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4639
  signal tmp_ivl_35395 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4639
  signal tmp_ivl_35400 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4639
  signal tmp_ivl_35403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4639
  signal tmp_ivl_35407 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4639
  signal tmp_ivl_35409 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4639
  signal tmp_ivl_3541 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3062
  signal tmp_ivl_35411 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4639
  signal tmp_ivl_35416 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4640
  signal tmp_ivl_3542 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3062
  signal tmp_ivl_35421 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4640
  signal tmp_ivl_35423 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4640
  signal tmp_ivl_35428 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4640
  signal tmp_ivl_35431 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4640
  signal tmp_ivl_35435 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4640
  signal tmp_ivl_35437 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4640
  signal tmp_ivl_35439 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4640
  signal tmp_ivl_35445 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4641
  signal tmp_ivl_35446 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4641
  signal tmp_ivl_35451 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4641
  signal tmp_ivl_35453 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4641
  signal tmp_ivl_35458 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4641
  signal tmp_ivl_35461 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4641
  signal tmp_ivl_35465 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4641
  signal tmp_ivl_35467 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4641
  signal tmp_ivl_35469 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4641
  signal tmp_ivl_3547 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3062
  signal tmp_ivl_35474 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4642
  signal tmp_ivl_35479 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4642
  signal tmp_ivl_35481 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4642
  signal tmp_ivl_35486 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4642
  signal tmp_ivl_35489 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4642
  signal tmp_ivl_35493 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4642
  signal tmp_ivl_35495 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4642
  signal tmp_ivl_35497 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4642
  signal tmp_ivl_3550 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3062
  signal tmp_ivl_35502 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4643
  signal tmp_ivl_35507 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4643
  signal tmp_ivl_35509 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4643
  signal tmp_ivl_35514 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4643
  signal tmp_ivl_35517 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4643
  signal tmp_ivl_3552 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3062
  signal tmp_ivl_35521 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4643
  signal tmp_ivl_35523 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4643
  signal tmp_ivl_35525 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4643
  signal tmp_ivl_3553 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3062
  signal tmp_ivl_35530 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4644
  signal tmp_ivl_35535 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4644
  signal tmp_ivl_35537 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4644
  signal tmp_ivl_35542 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4644
  signal tmp_ivl_35545 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4644
  signal tmp_ivl_35549 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4644
  signal tmp_ivl_35551 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4644
  signal tmp_ivl_35553 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4644
  signal tmp_ivl_35558 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4645
  signal tmp_ivl_35563 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4645
  signal tmp_ivl_35565 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4645
  signal tmp_ivl_35570 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4645
  signal tmp_ivl_35573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4645
  signal tmp_ivl_35577 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4645
  signal tmp_ivl_35579 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4645
  signal tmp_ivl_3558 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3062
  signal tmp_ivl_35581 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4645
  signal tmp_ivl_35586 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4646
  signal tmp_ivl_35591 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4646
  signal tmp_ivl_35593 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4646
  signal tmp_ivl_35598 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4646
  signal tmp_ivl_3560 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3062
  signal tmp_ivl_35601 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4646
  signal tmp_ivl_35605 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4646
  signal tmp_ivl_35607 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4646
  signal tmp_ivl_35609 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4646
  signal tmp_ivl_35614 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4647
  signal tmp_ivl_35619 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4647
  signal tmp_ivl_3562 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3062
  signal tmp_ivl_35621 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4647
  signal tmp_ivl_35626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4647
  signal tmp_ivl_35629 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4647
  signal tmp_ivl_35633 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4647
  signal tmp_ivl_35635 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4647
  signal tmp_ivl_35637 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4647
  signal tmp_ivl_35642 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4648
  signal tmp_ivl_35647 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4648
  signal tmp_ivl_35649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4648
  signal tmp_ivl_35654 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4648
  signal tmp_ivl_35657 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4648
  signal tmp_ivl_35661 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4648
  signal tmp_ivl_35663 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4648
  signal tmp_ivl_35665 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4648
  signal tmp_ivl_35670 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4649
  signal tmp_ivl_35675 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4649
  signal tmp_ivl_35677 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4649
  signal tmp_ivl_3568 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3063
  signal tmp_ivl_35682 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4649
  signal tmp_ivl_35685 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4649
  signal tmp_ivl_35689 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4649
  signal tmp_ivl_35691 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4649
  signal tmp_ivl_35693 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4649
  signal tmp_ivl_35698 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4650
  signal tmp_ivl_357 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2952
  signal tmp_ivl_3570 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3063
  signal tmp_ivl_35703 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4650
  signal tmp_ivl_35705 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4650
  signal tmp_ivl_3571 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3063
  signal tmp_ivl_35710 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4650
  signal tmp_ivl_35713 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4650
  signal tmp_ivl_35717 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4650
  signal tmp_ivl_35719 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4650
  signal tmp_ivl_35721 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4650
  signal tmp_ivl_35726 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4651
  signal tmp_ivl_35731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4651
  signal tmp_ivl_35733 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4651
  signal tmp_ivl_35738 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4651
  signal tmp_ivl_35741 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4651
  signal tmp_ivl_35745 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4651
  signal tmp_ivl_35747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4651
  signal tmp_ivl_35749 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4651
  signal tmp_ivl_35754 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4652
  signal tmp_ivl_35759 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4652
  signal tmp_ivl_3576 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3063
  signal tmp_ivl_35761 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4652
  signal tmp_ivl_35766 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4652
  signal tmp_ivl_35769 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4652
  signal tmp_ivl_35773 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4652
  signal tmp_ivl_35775 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4652
  signal tmp_ivl_35777 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4652
  signal tmp_ivl_35782 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4653
  signal tmp_ivl_35787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4653
  signal tmp_ivl_35789 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4653
  signal tmp_ivl_3579 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3063
  signal tmp_ivl_35794 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4653
  signal tmp_ivl_35797 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4653
  signal tmp_ivl_35801 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4653
  signal tmp_ivl_35803 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4653
  signal tmp_ivl_35805 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4653
  signal tmp_ivl_3581 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3063
  signal tmp_ivl_35810 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4654
  signal tmp_ivl_35815 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4654
  signal tmp_ivl_35817 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4654
  signal tmp_ivl_3582 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3063
  signal tmp_ivl_35822 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4654
  signal tmp_ivl_35825 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4654
  signal tmp_ivl_35829 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4654
  signal tmp_ivl_35831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4654
  signal tmp_ivl_35833 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4654
  signal tmp_ivl_35838 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4655
  signal tmp_ivl_35843 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4655
  signal tmp_ivl_35845 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4655
  signal tmp_ivl_35850 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4655
  signal tmp_ivl_35853 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4655
  signal tmp_ivl_35857 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4655
  signal tmp_ivl_35859 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4655
  signal tmp_ivl_35861 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4655
  signal tmp_ivl_35866 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4656
  signal tmp_ivl_3587 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3063
  signal tmp_ivl_35871 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4656
  signal tmp_ivl_35873 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4656
  signal tmp_ivl_35878 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4656
  signal tmp_ivl_35881 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4656
  signal tmp_ivl_35885 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4656
  signal tmp_ivl_35887 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4656
  signal tmp_ivl_35889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4656
  signal tmp_ivl_3589 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3063
  signal tmp_ivl_35894 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4657
  signal tmp_ivl_35899 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4657
  signal tmp_ivl_35901 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4657
  signal tmp_ivl_35906 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4657
  signal tmp_ivl_35909 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4657
  signal tmp_ivl_3591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3063
  signal tmp_ivl_35913 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4657
  signal tmp_ivl_35915 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4657
  signal tmp_ivl_35917 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4657
  signal tmp_ivl_35922 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4658
  signal tmp_ivl_35927 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4658
  signal tmp_ivl_35929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4658
  signal tmp_ivl_35934 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4658
  signal tmp_ivl_35937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4658
  signal tmp_ivl_35941 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4658
  signal tmp_ivl_35943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4658
  signal tmp_ivl_35945 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4658
  signal tmp_ivl_35950 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4659
  signal tmp_ivl_35955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4659
  signal tmp_ivl_35957 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4659
  signal tmp_ivl_35962 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4659
  signal tmp_ivl_35965 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4659
  signal tmp_ivl_35969 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4659
  signal tmp_ivl_3597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3064
  signal tmp_ivl_35971 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4659
  signal tmp_ivl_35973 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4659
  signal tmp_ivl_35978 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4660
  signal tmp_ivl_35983 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4660
  signal tmp_ivl_35985 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4660
  signal tmp_ivl_3599 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3064
  signal tmp_ivl_35990 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4660
  signal tmp_ivl_35993 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4660
  signal tmp_ivl_35997 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4660
  signal tmp_ivl_35999 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4660
  signal tmp_ivl_360 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2952
  signal tmp_ivl_3600 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3064
  signal tmp_ivl_36001 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4660
  signal tmp_ivl_36006 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4661
  signal tmp_ivl_36011 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4661
  signal tmp_ivl_36013 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4661
  signal tmp_ivl_36018 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4661
  signal tmp_ivl_36021 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4661
  signal tmp_ivl_36025 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4661
  signal tmp_ivl_36027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4661
  signal tmp_ivl_36029 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4661
  signal tmp_ivl_36034 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4662
  signal tmp_ivl_36039 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4662
  signal tmp_ivl_36041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4662
  signal tmp_ivl_36046 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4662
  signal tmp_ivl_36049 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4662
  signal tmp_ivl_3605 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3064
  signal tmp_ivl_36053 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4662
  signal tmp_ivl_36055 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4662
  signal tmp_ivl_36057 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4662
  signal tmp_ivl_36062 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4663
  signal tmp_ivl_36067 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4663
  signal tmp_ivl_36069 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4663
  signal tmp_ivl_36074 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4663
  signal tmp_ivl_36077 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4663
  signal tmp_ivl_3608 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3064
  signal tmp_ivl_36081 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4663
  signal tmp_ivl_36083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4663
  signal tmp_ivl_36085 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4663
  signal tmp_ivl_36090 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4664
  signal tmp_ivl_36095 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4664
  signal tmp_ivl_36097 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4664
  signal tmp_ivl_3610 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3064
  signal tmp_ivl_36102 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4664
  signal tmp_ivl_36105 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4664
  signal tmp_ivl_36109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4664
  signal tmp_ivl_3611 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3064
  signal tmp_ivl_36111 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4664
  signal tmp_ivl_36113 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4664
  signal tmp_ivl_36118 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4665
  signal tmp_ivl_36123 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4665
  signal tmp_ivl_36125 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4665
  signal tmp_ivl_36130 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4665
  signal tmp_ivl_36133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4665
  signal tmp_ivl_36137 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4665
  signal tmp_ivl_36139 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4665
  signal tmp_ivl_36141 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4665
  signal tmp_ivl_36146 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4666
  signal tmp_ivl_36151 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4666
  signal tmp_ivl_36153 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4666
  signal tmp_ivl_36158 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4666
  signal tmp_ivl_3616 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3064
  signal tmp_ivl_36161 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4666
  signal tmp_ivl_36165 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4666
  signal tmp_ivl_36167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4666
  signal tmp_ivl_36169 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4666
  signal tmp_ivl_36174 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4667
  signal tmp_ivl_36179 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4667
  signal tmp_ivl_3618 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3064
  signal tmp_ivl_36181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4667
  signal tmp_ivl_36186 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4667
  signal tmp_ivl_36189 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4667
  signal tmp_ivl_36193 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4667
  signal tmp_ivl_36195 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4667
  signal tmp_ivl_36197 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4667
  signal tmp_ivl_362 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2952
  signal tmp_ivl_3620 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3064
  signal tmp_ivl_36202 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4668
  signal tmp_ivl_36207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4668
  signal tmp_ivl_36209 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4668
  signal tmp_ivl_36214 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4668
  signal tmp_ivl_36217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4668
  signal tmp_ivl_36221 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4668
  signal tmp_ivl_36223 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4668
  signal tmp_ivl_36225 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4668
  signal tmp_ivl_36230 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4669
  signal tmp_ivl_36235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4669
  signal tmp_ivl_36237 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4669
  signal tmp_ivl_36242 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4669
  signal tmp_ivl_36245 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4669
  signal tmp_ivl_36249 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4669
  signal tmp_ivl_36251 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4669
  signal tmp_ivl_36253 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4669
  signal tmp_ivl_36258 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4670
  signal tmp_ivl_3626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3065
  signal tmp_ivl_36263 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4670
  signal tmp_ivl_36265 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4670
  signal tmp_ivl_36270 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4670
  signal tmp_ivl_36273 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4670
  signal tmp_ivl_36277 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4670
  signal tmp_ivl_36279 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4670
  signal tmp_ivl_3628 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3065
  signal tmp_ivl_36281 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4670
  signal tmp_ivl_36286 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4671
  signal tmp_ivl_3629 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3065
  signal tmp_ivl_36291 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4671
  signal tmp_ivl_36293 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4671
  signal tmp_ivl_36298 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4671
  signal tmp_ivl_363 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2952
  signal tmp_ivl_36301 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4671
  signal tmp_ivl_36305 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4671
  signal tmp_ivl_36307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4671
  signal tmp_ivl_36309 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4671
  signal tmp_ivl_36314 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4672
  signal tmp_ivl_36319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4672
  signal tmp_ivl_36321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4672
  signal tmp_ivl_36326 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4672
  signal tmp_ivl_36329 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4672
  signal tmp_ivl_36333 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4672
  signal tmp_ivl_36335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4672
  signal tmp_ivl_36337 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4672
  signal tmp_ivl_3634 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3065
  signal tmp_ivl_36342 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4673
  signal tmp_ivl_36347 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4673
  signal tmp_ivl_36349 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4673
  signal tmp_ivl_36354 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4673
  signal tmp_ivl_36357 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4673
  signal tmp_ivl_36361 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4673
  signal tmp_ivl_36363 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4673
  signal tmp_ivl_36365 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4673
  signal tmp_ivl_3637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3065
  signal tmp_ivl_36370 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4674
  signal tmp_ivl_36375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4674
  signal tmp_ivl_36377 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4674
  signal tmp_ivl_36382 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4674
  signal tmp_ivl_36385 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4674
  signal tmp_ivl_36389 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4674
  signal tmp_ivl_3639 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3065
  signal tmp_ivl_36391 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4674
  signal tmp_ivl_36393 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4674
  signal tmp_ivl_36398 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4675
  signal tmp_ivl_3640 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3065
  signal tmp_ivl_36403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4675
  signal tmp_ivl_36405 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4675
  signal tmp_ivl_36410 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4675
  signal tmp_ivl_36413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4675
  signal tmp_ivl_36417 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4675
  signal tmp_ivl_36419 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4675
  signal tmp_ivl_36421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4675
  signal tmp_ivl_36426 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4676
  signal tmp_ivl_36431 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4676
  signal tmp_ivl_36433 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4676
  signal tmp_ivl_36438 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4676
  signal tmp_ivl_36441 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4676
  signal tmp_ivl_36445 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4676
  signal tmp_ivl_36447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4676
  signal tmp_ivl_36449 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4676
  signal tmp_ivl_3645 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3065
  signal tmp_ivl_36454 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4677
  signal tmp_ivl_36459 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4677
  signal tmp_ivl_36461 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4677
  signal tmp_ivl_36466 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4677
  signal tmp_ivl_36469 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4677
  signal tmp_ivl_3647 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3065
  signal tmp_ivl_36473 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4677
  signal tmp_ivl_36475 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4677
  signal tmp_ivl_36477 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4677
  signal tmp_ivl_36482 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4678
  signal tmp_ivl_36487 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4678
  signal tmp_ivl_36489 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4678
  signal tmp_ivl_3649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3065
  signal tmp_ivl_36494 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4678
  signal tmp_ivl_36497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4678
  signal tmp_ivl_36501 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4678
  signal tmp_ivl_36503 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4678
  signal tmp_ivl_36505 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4678
  signal tmp_ivl_36510 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4679
  signal tmp_ivl_36515 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4679
  signal tmp_ivl_36517 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4679
  signal tmp_ivl_36522 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4679
  signal tmp_ivl_36525 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4679
  signal tmp_ivl_36529 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4679
  signal tmp_ivl_36531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4679
  signal tmp_ivl_36533 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4679
  signal tmp_ivl_36538 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4680
  signal tmp_ivl_36543 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4680
  signal tmp_ivl_36545 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4680
  signal tmp_ivl_3655 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3066
  signal tmp_ivl_36550 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4680
  signal tmp_ivl_36553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4680
  signal tmp_ivl_36557 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4680
  signal tmp_ivl_36559 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4680
  signal tmp_ivl_36561 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4680
  signal tmp_ivl_36566 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4681
  signal tmp_ivl_3657 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3066
  signal tmp_ivl_36571 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4681
  signal tmp_ivl_36573 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4681
  signal tmp_ivl_36578 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4681
  signal tmp_ivl_3658 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3066
  signal tmp_ivl_36581 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4681
  signal tmp_ivl_36585 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4681
  signal tmp_ivl_36587 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4681
  signal tmp_ivl_36589 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4681
  signal tmp_ivl_36594 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4682
  signal tmp_ivl_36599 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4682
  signal tmp_ivl_36601 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4682
  signal tmp_ivl_36606 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4682
  signal tmp_ivl_36609 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4682
  signal tmp_ivl_36613 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4682
  signal tmp_ivl_36615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4682
  signal tmp_ivl_36617 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4682
  signal tmp_ivl_36622 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4683
  signal tmp_ivl_36627 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4683
  signal tmp_ivl_36629 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4683
  signal tmp_ivl_3663 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3066
  signal tmp_ivl_36634 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4683
  signal tmp_ivl_36637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4683
  signal tmp_ivl_36641 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4683
  signal tmp_ivl_36643 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4683
  signal tmp_ivl_36645 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4683
  signal tmp_ivl_36650 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4684
  signal tmp_ivl_36655 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4684
  signal tmp_ivl_36657 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4684
  signal tmp_ivl_3666 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3066
  signal tmp_ivl_36662 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4684
  signal tmp_ivl_36665 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4684
  signal tmp_ivl_36669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4684
  signal tmp_ivl_36671 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4684
  signal tmp_ivl_36673 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4684
  signal tmp_ivl_36678 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4685
  signal tmp_ivl_3668 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3066
  signal tmp_ivl_36683 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4685
  signal tmp_ivl_36685 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4685
  signal tmp_ivl_3669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3066
  signal tmp_ivl_36690 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4685
  signal tmp_ivl_36693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4685
  signal tmp_ivl_36697 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4685
  signal tmp_ivl_36699 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4685
  signal tmp_ivl_36701 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4685
  signal tmp_ivl_36706 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4686
  signal tmp_ivl_36711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4686
  signal tmp_ivl_36713 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4686
  signal tmp_ivl_36718 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4686
  signal tmp_ivl_36721 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4686
  signal tmp_ivl_36725 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4686
  signal tmp_ivl_36727 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4686
  signal tmp_ivl_36729 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4686
  signal tmp_ivl_36734 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4687
  signal tmp_ivl_36739 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4687
  signal tmp_ivl_3674 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3066
  signal tmp_ivl_36741 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4687
  signal tmp_ivl_36746 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4687
  signal tmp_ivl_36749 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4687
  signal tmp_ivl_36753 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4687
  signal tmp_ivl_36755 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4687
  signal tmp_ivl_36757 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4687
  signal tmp_ivl_3676 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3066
  signal tmp_ivl_36762 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4688
  signal tmp_ivl_36767 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4688
  signal tmp_ivl_36769 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4688
  signal tmp_ivl_36774 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4688
  signal tmp_ivl_36777 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4688
  signal tmp_ivl_3678 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3066
  signal tmp_ivl_36781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4688
  signal tmp_ivl_36783 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4688
  signal tmp_ivl_36785 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4688
  signal tmp_ivl_36790 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4689
  signal tmp_ivl_36795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4689
  signal tmp_ivl_36797 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4689
  signal tmp_ivl_368 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2952
  signal tmp_ivl_36802 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4689
  signal tmp_ivl_36805 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4689
  signal tmp_ivl_36809 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4689
  signal tmp_ivl_36811 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4689
  signal tmp_ivl_36813 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4689
  signal tmp_ivl_36818 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4690
  signal tmp_ivl_36823 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4690
  signal tmp_ivl_36825 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4690
  signal tmp_ivl_36830 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4690
  signal tmp_ivl_36833 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4690
  signal tmp_ivl_36837 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4690
  signal tmp_ivl_36839 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4690
  signal tmp_ivl_3684 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3067
  signal tmp_ivl_36841 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4690
  signal tmp_ivl_36846 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4691
  signal tmp_ivl_36851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4691
  signal tmp_ivl_36853 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4691
  signal tmp_ivl_36858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4691
  signal tmp_ivl_3686 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3067
  signal tmp_ivl_36861 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4691
  signal tmp_ivl_36865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4691
  signal tmp_ivl_36867 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4691
  signal tmp_ivl_36869 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4691
  signal tmp_ivl_3687 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3067
  signal tmp_ivl_36874 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4692
  signal tmp_ivl_36879 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4692
  signal tmp_ivl_36881 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4692
  signal tmp_ivl_36886 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4692
  signal tmp_ivl_36889 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4692
  signal tmp_ivl_36893 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4692
  signal tmp_ivl_36895 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4692
  signal tmp_ivl_36897 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4692
  signal tmp_ivl_36902 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4693
  signal tmp_ivl_36907 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4693
  signal tmp_ivl_36909 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4693
  signal tmp_ivl_36914 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4693
  signal tmp_ivl_36917 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4693
  signal tmp_ivl_3692 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3067
  signal tmp_ivl_36921 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4693
  signal tmp_ivl_36923 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4693
  signal tmp_ivl_36925 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4693
  signal tmp_ivl_36931 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4694
  signal tmp_ivl_36932 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4694
  signal tmp_ivl_36937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4694
  signal tmp_ivl_36939 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4694
  signal tmp_ivl_36944 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4694
  signal tmp_ivl_36947 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4694
  signal tmp_ivl_3695 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3067
  signal tmp_ivl_36951 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4694
  signal tmp_ivl_36953 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4694
  signal tmp_ivl_36955 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4694
  signal tmp_ivl_36961 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4695
  signal tmp_ivl_36962 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4695
  signal tmp_ivl_36967 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4695
  signal tmp_ivl_36969 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4695
  signal tmp_ivl_3697 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3067
  signal tmp_ivl_36974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4695
  signal tmp_ivl_36977 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4695
  signal tmp_ivl_3698 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3067
  signal tmp_ivl_36981 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4695
  signal tmp_ivl_36983 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4695
  signal tmp_ivl_36985 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4695
  signal tmp_ivl_36991 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4696
  signal tmp_ivl_36992 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4696
  signal tmp_ivl_36997 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4696
  signal tmp_ivl_36999 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4696
  signal tmp_ivl_370 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2952
  signal tmp_ivl_37004 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4696
  signal tmp_ivl_37007 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4696
  signal tmp_ivl_37011 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4696
  signal tmp_ivl_37013 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4696
  signal tmp_ivl_37015 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4696
  signal tmp_ivl_37021 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4697
  signal tmp_ivl_37022 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4697
  signal tmp_ivl_37027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4697
  signal tmp_ivl_37029 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4697
  signal tmp_ivl_3703 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3067
  signal tmp_ivl_37034 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4697
  signal tmp_ivl_37037 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4697
  signal tmp_ivl_37041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4697
  signal tmp_ivl_37043 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4697
  signal tmp_ivl_37045 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4697
  signal tmp_ivl_3705 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3067
  signal tmp_ivl_37051 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4698
  signal tmp_ivl_37052 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4698
  signal tmp_ivl_37057 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4698
  signal tmp_ivl_37059 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4698
  signal tmp_ivl_37064 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4698
  signal tmp_ivl_37067 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4698
  signal tmp_ivl_3707 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3067
  signal tmp_ivl_37071 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4698
  signal tmp_ivl_37073 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4698
  signal tmp_ivl_37075 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4698
  signal tmp_ivl_37081 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4699
  signal tmp_ivl_37082 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4699
  signal tmp_ivl_37087 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4699
  signal tmp_ivl_37089 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4699
  signal tmp_ivl_37094 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4699
  signal tmp_ivl_37097 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4699
  signal tmp_ivl_37101 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4699
  signal tmp_ivl_37103 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4699
  signal tmp_ivl_37105 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4699
  signal tmp_ivl_37111 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4700
  signal tmp_ivl_37112 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4700
  signal tmp_ivl_37117 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4700
  signal tmp_ivl_37119 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4700
  signal tmp_ivl_37124 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4700
  signal tmp_ivl_37127 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4700
  signal tmp_ivl_3713 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3068
  signal tmp_ivl_37131 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4700
  signal tmp_ivl_37133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4700
  signal tmp_ivl_37135 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4700
  signal tmp_ivl_37141 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4701
  signal tmp_ivl_37142 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4701
  signal tmp_ivl_37147 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4701
  signal tmp_ivl_37149 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4701
  signal tmp_ivl_3715 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3068
  signal tmp_ivl_37154 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4701
  signal tmp_ivl_37157 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4701
  signal tmp_ivl_3716 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3068
  signal tmp_ivl_37161 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4701
  signal tmp_ivl_37163 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4701
  signal tmp_ivl_37165 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4701
  signal tmp_ivl_37171 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4702
  signal tmp_ivl_37172 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4702
  signal tmp_ivl_37177 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4702
  signal tmp_ivl_37179 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4702
  signal tmp_ivl_37184 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4702
  signal tmp_ivl_37187 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4702
  signal tmp_ivl_37191 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4702
  signal tmp_ivl_37193 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4702
  signal tmp_ivl_37195 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4702
  signal tmp_ivl_372 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2952
  signal tmp_ivl_37201 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4703
  signal tmp_ivl_37202 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4703
  signal tmp_ivl_37207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4703
  signal tmp_ivl_37209 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4703
  signal tmp_ivl_3721 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3068
  signal tmp_ivl_37214 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4703
  signal tmp_ivl_37217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4703
  signal tmp_ivl_37221 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4703
  signal tmp_ivl_37223 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4703
  signal tmp_ivl_37225 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4703
  signal tmp_ivl_37231 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4704
  signal tmp_ivl_37232 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4704
  signal tmp_ivl_37237 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4704
  signal tmp_ivl_37239 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4704
  signal tmp_ivl_3724 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3068
  signal tmp_ivl_37244 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4704
  signal tmp_ivl_37247 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4704
  signal tmp_ivl_37251 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4704
  signal tmp_ivl_37253 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4704
  signal tmp_ivl_37255 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4704
  signal tmp_ivl_3726 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3068
  signal tmp_ivl_37261 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4705
  signal tmp_ivl_37262 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4705
  signal tmp_ivl_37267 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4705
  signal tmp_ivl_37269 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4705
  signal tmp_ivl_3727 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3068
  signal tmp_ivl_37274 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4705
  signal tmp_ivl_37277 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4705
  signal tmp_ivl_37281 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4705
  signal tmp_ivl_37283 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4705
  signal tmp_ivl_37285 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4705
  signal tmp_ivl_37291 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4706
  signal tmp_ivl_37292 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4706
  signal tmp_ivl_37297 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4706
  signal tmp_ivl_37299 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4706
  signal tmp_ivl_37304 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4706
  signal tmp_ivl_37307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4706
  signal tmp_ivl_37311 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4706
  signal tmp_ivl_37313 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4706
  signal tmp_ivl_37315 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4706
  signal tmp_ivl_3732 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3068
  signal tmp_ivl_37321 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4707
  signal tmp_ivl_37322 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4707
  signal tmp_ivl_37327 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4707
  signal tmp_ivl_37329 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4707
  signal tmp_ivl_37334 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4707
  signal tmp_ivl_37337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4707
  signal tmp_ivl_3734 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3068
  signal tmp_ivl_37341 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4707
  signal tmp_ivl_37343 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4707
  signal tmp_ivl_37345 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4707
  signal tmp_ivl_37351 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4708
  signal tmp_ivl_37352 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4708
  signal tmp_ivl_37357 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4708
  signal tmp_ivl_37359 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4708
  signal tmp_ivl_37364 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4708
  signal tmp_ivl_37367 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4708
  signal tmp_ivl_37371 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4708
  signal tmp_ivl_37373 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4708
  signal tmp_ivl_37375 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4708
  signal tmp_ivl_37381 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4709
  signal tmp_ivl_37382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4709
  signal tmp_ivl_37387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4709
  signal tmp_ivl_37389 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4709
  signal tmp_ivl_37394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4709
  signal tmp_ivl_37397 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4709
  signal tmp_ivl_3740 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3069
  signal tmp_ivl_37401 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4709
  signal tmp_ivl_37403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4709
  signal tmp_ivl_37405 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4709
  signal tmp_ivl_37411 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4710
  signal tmp_ivl_37412 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4710
  signal tmp_ivl_37417 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4710
  signal tmp_ivl_37419 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4710
  signal tmp_ivl_3742 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3069
  signal tmp_ivl_37424 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4710
  signal tmp_ivl_37427 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4710
  signal tmp_ivl_3743 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3069
  signal tmp_ivl_37431 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4710
  signal tmp_ivl_37433 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4710
  signal tmp_ivl_37435 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4710
  signal tmp_ivl_37441 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4711
  signal tmp_ivl_37442 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4711
  signal tmp_ivl_37447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4711
  signal tmp_ivl_37449 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4711
  signal tmp_ivl_37454 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4711
  signal tmp_ivl_37457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4711
  signal tmp_ivl_37461 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4711
  signal tmp_ivl_37463 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4711
  signal tmp_ivl_37465 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4711
  signal tmp_ivl_37471 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4712
  signal tmp_ivl_37472 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4712
  signal tmp_ivl_37477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4712
  signal tmp_ivl_37479 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4712
  signal tmp_ivl_3748 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3069
  signal tmp_ivl_37484 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4712
  signal tmp_ivl_37487 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4712
  signal tmp_ivl_37491 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4712
  signal tmp_ivl_37493 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4712
  signal tmp_ivl_37495 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4712
  signal tmp_ivl_37501 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4713
  signal tmp_ivl_37502 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4713
  signal tmp_ivl_37507 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4713
  signal tmp_ivl_37509 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4713
  signal tmp_ivl_3751 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3069
  signal tmp_ivl_37514 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4713
  signal tmp_ivl_37517 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4713
  signal tmp_ivl_37521 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4713
  signal tmp_ivl_37523 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4713
  signal tmp_ivl_37525 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4713
  signal tmp_ivl_3753 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3069
  signal tmp_ivl_37531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4714
  signal tmp_ivl_37532 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4714
  signal tmp_ivl_37537 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4714
  signal tmp_ivl_37539 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4714
  signal tmp_ivl_3754 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3069
  signal tmp_ivl_37544 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4714
  signal tmp_ivl_37547 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4714
  signal tmp_ivl_37551 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4714
  signal tmp_ivl_37553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4714
  signal tmp_ivl_37555 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4714
  signal tmp_ivl_37561 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4715
  signal tmp_ivl_37562 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4715
  signal tmp_ivl_37567 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4715
  signal tmp_ivl_37569 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4715
  signal tmp_ivl_37574 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4715
  signal tmp_ivl_37577 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4715
  signal tmp_ivl_37581 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4715
  signal tmp_ivl_37583 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4715
  signal tmp_ivl_37585 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4715
  signal tmp_ivl_3759 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3069
  signal tmp_ivl_37591 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4716
  signal tmp_ivl_37592 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4716
  signal tmp_ivl_37597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4716
  signal tmp_ivl_37599 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4716
  signal tmp_ivl_37604 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4716
  signal tmp_ivl_37607 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4716
  signal tmp_ivl_3761 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3069
  signal tmp_ivl_37611 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4716
  signal tmp_ivl_37613 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4716
  signal tmp_ivl_37615 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4716
  signal tmp_ivl_37621 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4717
  signal tmp_ivl_37622 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4717
  signal tmp_ivl_37627 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4717
  signal tmp_ivl_37629 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4717
  signal tmp_ivl_37634 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4717
  signal tmp_ivl_37637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4717
  signal tmp_ivl_37641 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4717
  signal tmp_ivl_37643 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4717
  signal tmp_ivl_37645 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4717
  signal tmp_ivl_37651 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4718
  signal tmp_ivl_37652 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4718
  signal tmp_ivl_37657 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4718
  signal tmp_ivl_37659 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4718
  signal tmp_ivl_37664 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4718
  signal tmp_ivl_37667 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4718
  signal tmp_ivl_3767 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3070
  signal tmp_ivl_37671 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4718
  signal tmp_ivl_37673 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4718
  signal tmp_ivl_37675 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4718
  signal tmp_ivl_37681 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4719
  signal tmp_ivl_37682 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4719
  signal tmp_ivl_37687 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4719
  signal tmp_ivl_37689 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4719
  signal tmp_ivl_3769 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3070
  signal tmp_ivl_37694 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4719
  signal tmp_ivl_37697 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4719
  signal tmp_ivl_3770 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3070
  signal tmp_ivl_37701 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4719
  signal tmp_ivl_37703 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4719
  signal tmp_ivl_37705 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4719
  signal tmp_ivl_37711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4720
  signal tmp_ivl_37712 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4720
  signal tmp_ivl_37717 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4720
  signal tmp_ivl_37719 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4720
  signal tmp_ivl_37724 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4720
  signal tmp_ivl_37727 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4720
  signal tmp_ivl_37731 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4720
  signal tmp_ivl_37733 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4720
  signal tmp_ivl_37735 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4720
  signal tmp_ivl_37741 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4721
  signal tmp_ivl_37742 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4721
  signal tmp_ivl_37747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4721
  signal tmp_ivl_37749 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4721
  signal tmp_ivl_3775 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3070
  signal tmp_ivl_37754 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4721
  signal tmp_ivl_37757 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4721
  signal tmp_ivl_37761 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4721
  signal tmp_ivl_37763 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4721
  signal tmp_ivl_37765 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4721
  signal tmp_ivl_37771 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4722
  signal tmp_ivl_37772 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4722
  signal tmp_ivl_37777 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4722
  signal tmp_ivl_37779 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4722
  signal tmp_ivl_3778 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3070
  signal tmp_ivl_37784 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4722
  signal tmp_ivl_37787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4722
  signal tmp_ivl_37791 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4722
  signal tmp_ivl_37793 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4722
  signal tmp_ivl_37795 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4722
  signal tmp_ivl_378 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2953
  signal tmp_ivl_3780 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3070
  signal tmp_ivl_37801 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4723
  signal tmp_ivl_37802 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4723
  signal tmp_ivl_37807 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4723
  signal tmp_ivl_37809 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4723
  signal tmp_ivl_3781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3070
  signal tmp_ivl_37814 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4723
  signal tmp_ivl_37817 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4723
  signal tmp_ivl_37821 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4723
  signal tmp_ivl_37823 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4723
  signal tmp_ivl_37825 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4723
  signal tmp_ivl_37831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4724
  signal tmp_ivl_37832 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4724
  signal tmp_ivl_37837 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4724
  signal tmp_ivl_37839 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4724
  signal tmp_ivl_37844 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4724
  signal tmp_ivl_37847 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4724
  signal tmp_ivl_37851 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4724
  signal tmp_ivl_37853 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4724
  signal tmp_ivl_37855 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4724
  signal tmp_ivl_3786 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3070
  signal tmp_ivl_37861 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4725
  signal tmp_ivl_37862 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4725
  signal tmp_ivl_37867 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4725
  signal tmp_ivl_37869 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4725
  signal tmp_ivl_37874 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4725
  signal tmp_ivl_37877 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4725
  signal tmp_ivl_3788 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3070
  signal tmp_ivl_37881 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4725
  signal tmp_ivl_37883 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4725
  signal tmp_ivl_37885 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4725
  signal tmp_ivl_37891 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4726
  signal tmp_ivl_37892 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4726
  signal tmp_ivl_37897 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4726
  signal tmp_ivl_37899 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4726
  signal tmp_ivl_37904 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4726
  signal tmp_ivl_37907 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4726
  signal tmp_ivl_37911 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4726
  signal tmp_ivl_37913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4726
  signal tmp_ivl_37915 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4726
  signal tmp_ivl_37921 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4727
  signal tmp_ivl_37922 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4727
  signal tmp_ivl_37927 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4727
  signal tmp_ivl_37929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4727
  signal tmp_ivl_37934 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4727
  signal tmp_ivl_37937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4727
  signal tmp_ivl_3794 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3071
  signal tmp_ivl_37941 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4727
  signal tmp_ivl_37943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4727
  signal tmp_ivl_37945 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4727
  signal tmp_ivl_37951 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4728
  signal tmp_ivl_37952 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4728
  signal tmp_ivl_37957 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4728
  signal tmp_ivl_37959 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4728
  signal tmp_ivl_3796 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3071
  signal tmp_ivl_37964 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4728
  signal tmp_ivl_37967 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4728
  signal tmp_ivl_3797 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3071
  signal tmp_ivl_37971 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4728
  signal tmp_ivl_37973 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4728
  signal tmp_ivl_37975 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4728
  signal tmp_ivl_37981 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4729
  signal tmp_ivl_37982 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4729
  signal tmp_ivl_37987 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4729
  signal tmp_ivl_37989 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4729
  signal tmp_ivl_37994 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4729
  signal tmp_ivl_37997 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4729
  signal tmp_ivl_38 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2941
  signal tmp_ivl_380 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2953
  signal tmp_ivl_38001 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4729
  signal tmp_ivl_38003 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4729
  signal tmp_ivl_38005 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4729
  signal tmp_ivl_38011 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4730
  signal tmp_ivl_38012 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4730
  signal tmp_ivl_38017 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4730
  signal tmp_ivl_38019 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4730
  signal tmp_ivl_3802 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3071
  signal tmp_ivl_38024 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4730
  signal tmp_ivl_38027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4730
  signal tmp_ivl_38031 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4730
  signal tmp_ivl_38033 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4730
  signal tmp_ivl_38035 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4730
  signal tmp_ivl_38041 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4731
  signal tmp_ivl_38042 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4731
  signal tmp_ivl_38047 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4731
  signal tmp_ivl_38049 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4731
  signal tmp_ivl_3805 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3071
  signal tmp_ivl_38054 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4731
  signal tmp_ivl_38057 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4731
  signal tmp_ivl_38061 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4731
  signal tmp_ivl_38063 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4731
  signal tmp_ivl_38065 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4731
  signal tmp_ivl_3807 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3071
  signal tmp_ivl_38071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4732
  signal tmp_ivl_38072 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4732
  signal tmp_ivl_38077 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4732
  signal tmp_ivl_38079 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4732
  signal tmp_ivl_3808 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3071
  signal tmp_ivl_38084 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4732
  signal tmp_ivl_38087 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4732
  signal tmp_ivl_38091 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4732
  signal tmp_ivl_38093 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4732
  signal tmp_ivl_38095 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4732
  signal tmp_ivl_381 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2953
  signal tmp_ivl_38101 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4733
  signal tmp_ivl_38102 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4733
  signal tmp_ivl_38107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4733
  signal tmp_ivl_38109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4733
  signal tmp_ivl_38114 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4733
  signal tmp_ivl_38117 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4733
  signal tmp_ivl_38121 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4733
  signal tmp_ivl_38123 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4733
  signal tmp_ivl_38125 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4733
  signal tmp_ivl_3813 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3071
  signal tmp_ivl_38131 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4734
  signal tmp_ivl_38132 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4734
  signal tmp_ivl_38137 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4734
  signal tmp_ivl_38139 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4734
  signal tmp_ivl_38144 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4734
  signal tmp_ivl_38147 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4734
  signal tmp_ivl_3815 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3071
  signal tmp_ivl_38151 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4734
  signal tmp_ivl_38153 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4734
  signal tmp_ivl_38155 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4734
  signal tmp_ivl_38161 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4735
  signal tmp_ivl_38162 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4735
  signal tmp_ivl_38167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4735
  signal tmp_ivl_38169 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4735
  signal tmp_ivl_38174 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4735
  signal tmp_ivl_38177 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4735
  signal tmp_ivl_38181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4735
  signal tmp_ivl_38183 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4735
  signal tmp_ivl_38185 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4735
  signal tmp_ivl_38191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4736
  signal tmp_ivl_38192 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4736
  signal tmp_ivl_38197 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4736
  signal tmp_ivl_38199 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4736
  signal tmp_ivl_38204 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4736
  signal tmp_ivl_38207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4736
  signal tmp_ivl_3821 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3072
  signal tmp_ivl_38211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4736
  signal tmp_ivl_38213 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4736
  signal tmp_ivl_38215 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4736
  signal tmp_ivl_38221 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4737
  signal tmp_ivl_38222 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4737
  signal tmp_ivl_38227 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4737
  signal tmp_ivl_38229 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4737
  signal tmp_ivl_3823 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3072
  signal tmp_ivl_38234 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4737
  signal tmp_ivl_38237 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4737
  signal tmp_ivl_3824 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3072
  signal tmp_ivl_38241 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4737
  signal tmp_ivl_38243 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4737
  signal tmp_ivl_38245 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4737
  signal tmp_ivl_38251 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4738
  signal tmp_ivl_38252 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4738
  signal tmp_ivl_38257 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4738
  signal tmp_ivl_38259 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4738
  signal tmp_ivl_38264 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4738
  signal tmp_ivl_38267 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4738
  signal tmp_ivl_38271 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4738
  signal tmp_ivl_38273 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4738
  signal tmp_ivl_38275 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4738
  signal tmp_ivl_38281 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4739
  signal tmp_ivl_38282 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4739
  signal tmp_ivl_38287 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4739
  signal tmp_ivl_38289 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4739
  signal tmp_ivl_3829 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3072
  signal tmp_ivl_38294 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4739
  signal tmp_ivl_38297 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4739
  signal tmp_ivl_38301 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4739
  signal tmp_ivl_38303 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4739
  signal tmp_ivl_38305 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4739
  signal tmp_ivl_38311 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4740
  signal tmp_ivl_38312 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4740
  signal tmp_ivl_38317 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4740
  signal tmp_ivl_38319 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4740
  signal tmp_ivl_3832 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3072
  signal tmp_ivl_38324 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4740
  signal tmp_ivl_38327 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4740
  signal tmp_ivl_38331 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4740
  signal tmp_ivl_38333 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4740
  signal tmp_ivl_38335 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4740
  signal tmp_ivl_3834 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3072
  signal tmp_ivl_38341 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4741
  signal tmp_ivl_38342 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4741
  signal tmp_ivl_38347 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4741
  signal tmp_ivl_38349 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4741
  signal tmp_ivl_3835 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3072
  signal tmp_ivl_38354 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4741
  signal tmp_ivl_38357 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4741
  signal tmp_ivl_38361 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4741
  signal tmp_ivl_38363 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4741
  signal tmp_ivl_38365 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4741
  signal tmp_ivl_38371 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4742
  signal tmp_ivl_38372 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4742
  signal tmp_ivl_38377 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4742
  signal tmp_ivl_38379 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4742
  signal tmp_ivl_38384 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4742
  signal tmp_ivl_38387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4742
  signal tmp_ivl_38391 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4742
  signal tmp_ivl_38393 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4742
  signal tmp_ivl_38395 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4742
  signal tmp_ivl_3840 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3072
  signal tmp_ivl_38401 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4743
  signal tmp_ivl_38402 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4743
  signal tmp_ivl_38407 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4743
  signal tmp_ivl_38409 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4743
  signal tmp_ivl_38414 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4743
  signal tmp_ivl_38417 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4743
  signal tmp_ivl_3842 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3072
  signal tmp_ivl_38421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4743
  signal tmp_ivl_38423 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4743
  signal tmp_ivl_38425 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4743
  signal tmp_ivl_38431 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4744
  signal tmp_ivl_38432 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4744
  signal tmp_ivl_38437 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4744
  signal tmp_ivl_38439 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4744
  signal tmp_ivl_38444 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4744
  signal tmp_ivl_38447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4744
  signal tmp_ivl_38451 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4744
  signal tmp_ivl_38453 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4744
  signal tmp_ivl_38455 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4744
  signal tmp_ivl_38461 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4745
  signal tmp_ivl_38462 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4745
  signal tmp_ivl_38467 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4745
  signal tmp_ivl_38469 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4745
  signal tmp_ivl_38474 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4745
  signal tmp_ivl_38477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4745
  signal tmp_ivl_3848 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3073
  signal tmp_ivl_38481 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4745
  signal tmp_ivl_38483 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4745
  signal tmp_ivl_38485 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4745
  signal tmp_ivl_38491 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4746
  signal tmp_ivl_38492 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4746
  signal tmp_ivl_38497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4746
  signal tmp_ivl_38499 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4746
  signal tmp_ivl_3850 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3073
  signal tmp_ivl_38504 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4746
  signal tmp_ivl_38507 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4746
  signal tmp_ivl_3851 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3073
  signal tmp_ivl_38511 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4746
  signal tmp_ivl_38513 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4746
  signal tmp_ivl_38515 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4746
  signal tmp_ivl_38521 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4747
  signal tmp_ivl_38522 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4747
  signal tmp_ivl_38527 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4747
  signal tmp_ivl_38529 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4747
  signal tmp_ivl_38534 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4747
  signal tmp_ivl_38537 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4747
  signal tmp_ivl_38541 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4747
  signal tmp_ivl_38543 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4747
  signal tmp_ivl_38545 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4747
  signal tmp_ivl_38551 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4748
  signal tmp_ivl_38552 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4748
  signal tmp_ivl_38557 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4748
  signal tmp_ivl_38559 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4748
  signal tmp_ivl_3856 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3073
  signal tmp_ivl_38564 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4748
  signal tmp_ivl_38567 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4748
  signal tmp_ivl_38571 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4748
  signal tmp_ivl_38573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4748
  signal tmp_ivl_38575 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4748
  signal tmp_ivl_38581 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4749
  signal tmp_ivl_38582 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4749
  signal tmp_ivl_38587 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4749
  signal tmp_ivl_38589 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4749
  signal tmp_ivl_3859 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3073
  signal tmp_ivl_38594 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4749
  signal tmp_ivl_38597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4749
  signal tmp_ivl_386 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2953
  signal tmp_ivl_38601 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4749
  signal tmp_ivl_38603 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4749
  signal tmp_ivl_38605 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4749
  signal tmp_ivl_3861 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3073
  signal tmp_ivl_38611 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4750
  signal tmp_ivl_38612 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4750
  signal tmp_ivl_38617 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4750
  signal tmp_ivl_38619 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4750
  signal tmp_ivl_3862 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3073
  signal tmp_ivl_38624 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4750
  signal tmp_ivl_38627 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4750
  signal tmp_ivl_38631 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4750
  signal tmp_ivl_38633 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4750
  signal tmp_ivl_38635 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4750
  signal tmp_ivl_38641 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4751
  signal tmp_ivl_38642 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4751
  signal tmp_ivl_38647 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4751
  signal tmp_ivl_38649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4751
  signal tmp_ivl_38654 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4751
  signal tmp_ivl_38657 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4751
  signal tmp_ivl_38661 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4751
  signal tmp_ivl_38663 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4751
  signal tmp_ivl_38665 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4751
  signal tmp_ivl_3867 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3073
  signal tmp_ivl_38671 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4752
  signal tmp_ivl_38672 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4752
  signal tmp_ivl_38677 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4752
  signal tmp_ivl_38679 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4752
  signal tmp_ivl_38684 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4752
  signal tmp_ivl_38687 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4752
  signal tmp_ivl_3869 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3073
  signal tmp_ivl_38691 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4752
  signal tmp_ivl_38693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4752
  signal tmp_ivl_38695 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4752
  signal tmp_ivl_38701 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4753
  signal tmp_ivl_38702 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4753
  signal tmp_ivl_38707 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4753
  signal tmp_ivl_38709 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4753
  signal tmp_ivl_38714 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4753
  signal tmp_ivl_38717 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4753
  signal tmp_ivl_38721 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4753
  signal tmp_ivl_38723 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4753
  signal tmp_ivl_38725 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4753
  signal tmp_ivl_38731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4754
  signal tmp_ivl_38732 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4754
  signal tmp_ivl_38737 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4754
  signal tmp_ivl_38739 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4754
  signal tmp_ivl_38744 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4754
  signal tmp_ivl_38747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4754
  signal tmp_ivl_3875 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3074
  signal tmp_ivl_38751 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4754
  signal tmp_ivl_38753 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4754
  signal tmp_ivl_38755 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4754
  signal tmp_ivl_38761 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4755
  signal tmp_ivl_38762 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4755
  signal tmp_ivl_38767 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4755
  signal tmp_ivl_38769 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4755
  signal tmp_ivl_3877 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3074
  signal tmp_ivl_38774 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4755
  signal tmp_ivl_38777 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4755
  signal tmp_ivl_3878 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3074
  signal tmp_ivl_38781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4755
  signal tmp_ivl_38783 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4755
  signal tmp_ivl_38785 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4755
  signal tmp_ivl_38791 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4756
  signal tmp_ivl_38792 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4756
  signal tmp_ivl_38797 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4756
  signal tmp_ivl_38799 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4756
  signal tmp_ivl_38804 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4756
  signal tmp_ivl_38807 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4756
  signal tmp_ivl_38811 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4756
  signal tmp_ivl_38813 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4756
  signal tmp_ivl_38815 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4756
  signal tmp_ivl_38821 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4757
  signal tmp_ivl_38822 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4757
  signal tmp_ivl_38827 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4757
  signal tmp_ivl_38829 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4757
  signal tmp_ivl_3883 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3074
  signal tmp_ivl_38834 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4757
  signal tmp_ivl_38837 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4757
  signal tmp_ivl_38841 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4757
  signal tmp_ivl_38843 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4757
  signal tmp_ivl_38845 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4757
  signal tmp_ivl_38851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4758
  signal tmp_ivl_38852 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4758
  signal tmp_ivl_38857 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4758
  signal tmp_ivl_38859 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4758
  signal tmp_ivl_3886 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3074
  signal tmp_ivl_38864 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4758
  signal tmp_ivl_38867 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4758
  signal tmp_ivl_38871 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4758
  signal tmp_ivl_38873 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4758
  signal tmp_ivl_38875 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4758
  signal tmp_ivl_3888 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3074
  signal tmp_ivl_38881 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4759
  signal tmp_ivl_38882 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4759
  signal tmp_ivl_38887 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4759
  signal tmp_ivl_38889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4759
  signal tmp_ivl_3889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3074
  signal tmp_ivl_38894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4759
  signal tmp_ivl_38897 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4759
  signal tmp_ivl_389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2953
  signal tmp_ivl_38901 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4759
  signal tmp_ivl_38903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4759
  signal tmp_ivl_38905 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4759
  signal tmp_ivl_38911 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4760
  signal tmp_ivl_38912 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4760
  signal tmp_ivl_38917 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4760
  signal tmp_ivl_38919 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4760
  signal tmp_ivl_38924 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4760
  signal tmp_ivl_38927 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4760
  signal tmp_ivl_38931 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4760
  signal tmp_ivl_38933 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4760
  signal tmp_ivl_38935 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4760
  signal tmp_ivl_3894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3074
  signal tmp_ivl_38941 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4761
  signal tmp_ivl_38942 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4761
  signal tmp_ivl_38947 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4761
  signal tmp_ivl_38949 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4761
  signal tmp_ivl_38954 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4761
  signal tmp_ivl_38957 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4761
  signal tmp_ivl_3896 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3074
  signal tmp_ivl_38961 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4761
  signal tmp_ivl_38963 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4761
  signal tmp_ivl_38965 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4761
  signal tmp_ivl_38971 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4762
  signal tmp_ivl_38972 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4762
  signal tmp_ivl_38977 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4762
  signal tmp_ivl_38979 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4762
  signal tmp_ivl_38984 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4762
  signal tmp_ivl_38987 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4762
  signal tmp_ivl_38991 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4762
  signal tmp_ivl_38993 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4762
  signal tmp_ivl_38995 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4762
  signal tmp_ivl_39001 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4763
  signal tmp_ivl_39002 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4763
  signal tmp_ivl_39007 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4763
  signal tmp_ivl_39009 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4763
  signal tmp_ivl_39014 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4763
  signal tmp_ivl_39017 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4763
  signal tmp_ivl_3902 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3075
  signal tmp_ivl_39021 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4763
  signal tmp_ivl_39023 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4763
  signal tmp_ivl_39025 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4763
  signal tmp_ivl_39031 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4764
  signal tmp_ivl_39032 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4764
  signal tmp_ivl_39037 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4764
  signal tmp_ivl_39039 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4764
  signal tmp_ivl_3904 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3075
  signal tmp_ivl_39044 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4764
  signal tmp_ivl_39047 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4764
  signal tmp_ivl_3905 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3075
  signal tmp_ivl_39051 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4764
  signal tmp_ivl_39053 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4764
  signal tmp_ivl_39055 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4764
  signal tmp_ivl_39061 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4765
  signal tmp_ivl_39062 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4765
  signal tmp_ivl_39067 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4765
  signal tmp_ivl_39069 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4765
  signal tmp_ivl_39074 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4765
  signal tmp_ivl_39077 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4765
  signal tmp_ivl_39081 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4765
  signal tmp_ivl_39083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4765
  signal tmp_ivl_39085 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4765
  signal tmp_ivl_39091 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4766
  signal tmp_ivl_39092 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4766
  signal tmp_ivl_39097 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4766
  signal tmp_ivl_39099 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4766
  signal tmp_ivl_391 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2953
  signal tmp_ivl_3910 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3075
  signal tmp_ivl_39104 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4766
  signal tmp_ivl_39107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4766
  signal tmp_ivl_39111 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4766
  signal tmp_ivl_39113 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4766
  signal tmp_ivl_39115 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4766
  signal tmp_ivl_39121 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4767
  signal tmp_ivl_39122 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4767
  signal tmp_ivl_39127 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4767
  signal tmp_ivl_39129 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4767
  signal tmp_ivl_3913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3075
  signal tmp_ivl_39134 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4767
  signal tmp_ivl_39137 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4767
  signal tmp_ivl_39141 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4767
  signal tmp_ivl_39143 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4767
  signal tmp_ivl_39145 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4767
  signal tmp_ivl_3915 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3075
  signal tmp_ivl_39151 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4768
  signal tmp_ivl_39152 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4768
  signal tmp_ivl_39157 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4768
  signal tmp_ivl_39159 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4768
  signal tmp_ivl_3916 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3075
  signal tmp_ivl_39164 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4768
  signal tmp_ivl_39167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4768
  signal tmp_ivl_39171 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4768
  signal tmp_ivl_39173 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4768
  signal tmp_ivl_39175 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4768
  signal tmp_ivl_39181 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4769
  signal tmp_ivl_39182 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4769
  signal tmp_ivl_39187 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4769
  signal tmp_ivl_39189 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4769
  signal tmp_ivl_39194 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4769
  signal tmp_ivl_39197 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4769
  signal tmp_ivl_392 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2953
  signal tmp_ivl_39201 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4769
  signal tmp_ivl_39203 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4769
  signal tmp_ivl_39205 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4769
  signal tmp_ivl_3921 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3075
  signal tmp_ivl_39211 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4770
  signal tmp_ivl_39212 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4770
  signal tmp_ivl_39217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4770
  signal tmp_ivl_39219 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4770
  signal tmp_ivl_39224 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4770
  signal tmp_ivl_39227 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4770
  signal tmp_ivl_3923 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3075
  signal tmp_ivl_39231 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4770
  signal tmp_ivl_39233 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4770
  signal tmp_ivl_39235 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4770
  signal tmp_ivl_39241 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4771
  signal tmp_ivl_39242 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4771
  signal tmp_ivl_39247 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4771
  signal tmp_ivl_39249 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4771
  signal tmp_ivl_39254 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4771
  signal tmp_ivl_39257 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4771
  signal tmp_ivl_39261 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4771
  signal tmp_ivl_39263 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4771
  signal tmp_ivl_39265 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4771
  signal tmp_ivl_39271 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4772
  signal tmp_ivl_39272 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4772
  signal tmp_ivl_39277 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4772
  signal tmp_ivl_39279 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4772
  signal tmp_ivl_39284 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4772
  signal tmp_ivl_39287 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4772
  signal tmp_ivl_3929 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3076
  signal tmp_ivl_39291 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4772
  signal tmp_ivl_39293 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4772
  signal tmp_ivl_39295 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4772
  signal tmp_ivl_39301 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4773
  signal tmp_ivl_39302 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4773
  signal tmp_ivl_39307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4773
  signal tmp_ivl_39309 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4773
  signal tmp_ivl_3931 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3076
  signal tmp_ivl_39314 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4773
  signal tmp_ivl_39317 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4773
  signal tmp_ivl_3932 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3076
  signal tmp_ivl_39321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4773
  signal tmp_ivl_39323 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4773
  signal tmp_ivl_39325 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4773
  signal tmp_ivl_39331 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4774
  signal tmp_ivl_39332 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4774
  signal tmp_ivl_39337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4774
  signal tmp_ivl_39339 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4774
  signal tmp_ivl_39344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4774
  signal tmp_ivl_39347 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4774
  signal tmp_ivl_39351 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4774
  signal tmp_ivl_39353 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4774
  signal tmp_ivl_39355 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4774
  signal tmp_ivl_39361 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4775
  signal tmp_ivl_39362 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4775
  signal tmp_ivl_39367 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4775
  signal tmp_ivl_39369 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4775
  signal tmp_ivl_3937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3076
  signal tmp_ivl_39374 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4775
  signal tmp_ivl_39377 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4775
  signal tmp_ivl_39381 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4775
  signal tmp_ivl_39383 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4775
  signal tmp_ivl_39385 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4775
  signal tmp_ivl_39391 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4776
  signal tmp_ivl_39392 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4776
  signal tmp_ivl_39397 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4776
  signal tmp_ivl_39399 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4776
  signal tmp_ivl_3940 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3076
  signal tmp_ivl_39404 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4776
  signal tmp_ivl_39407 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4776
  signal tmp_ivl_39411 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4776
  signal tmp_ivl_39413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4776
  signal tmp_ivl_39415 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4776
  signal tmp_ivl_3942 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3076
  signal tmp_ivl_39421 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4777
  signal tmp_ivl_39422 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4777
  signal tmp_ivl_39427 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4777
  signal tmp_ivl_39429 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4777
  signal tmp_ivl_3943 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3076
  signal tmp_ivl_39434 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4777
  signal tmp_ivl_39437 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4777
  signal tmp_ivl_39441 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4777
  signal tmp_ivl_39443 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4777
  signal tmp_ivl_39445 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4777
  signal tmp_ivl_39451 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4778
  signal tmp_ivl_39452 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4778
  signal tmp_ivl_39457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4778
  signal tmp_ivl_39459 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4778
  signal tmp_ivl_39464 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4778
  signal tmp_ivl_39467 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4778
  signal tmp_ivl_39471 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4778
  signal tmp_ivl_39473 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4778
  signal tmp_ivl_39475 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4778
  signal tmp_ivl_3948 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3076
  signal tmp_ivl_39481 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4779
  signal tmp_ivl_39482 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4779
  signal tmp_ivl_39487 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4779
  signal tmp_ivl_39489 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4779
  signal tmp_ivl_39494 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4779
  signal tmp_ivl_39497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4779
  signal tmp_ivl_3950 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3076
  signal tmp_ivl_39501 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4779
  signal tmp_ivl_39503 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4779
  signal tmp_ivl_39505 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4779
  signal tmp_ivl_39511 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4780
  signal tmp_ivl_39512 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4780
  signal tmp_ivl_39517 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4780
  signal tmp_ivl_39519 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4780
  signal tmp_ivl_39524 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4780
  signal tmp_ivl_39527 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4780
  signal tmp_ivl_39531 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4780
  signal tmp_ivl_39533 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4780
  signal tmp_ivl_39535 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4780
  signal tmp_ivl_39541 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4781
  signal tmp_ivl_39542 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4781
  signal tmp_ivl_39547 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4781
  signal tmp_ivl_39549 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4781
  signal tmp_ivl_39554 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4781
  signal tmp_ivl_39557 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4781
  signal tmp_ivl_3956 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3077
  signal tmp_ivl_39561 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4781
  signal tmp_ivl_39563 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4781
  signal tmp_ivl_39565 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4781
  signal tmp_ivl_39571 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4782
  signal tmp_ivl_39572 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4782
  signal tmp_ivl_39577 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4782
  signal tmp_ivl_39579 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4782
  signal tmp_ivl_3958 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3077
  signal tmp_ivl_39584 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4782
  signal tmp_ivl_39587 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4782
  signal tmp_ivl_3959 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3077
  signal tmp_ivl_39591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4782
  signal tmp_ivl_39593 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4782
  signal tmp_ivl_39595 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4782
  signal tmp_ivl_39601 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4783
  signal tmp_ivl_39602 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4783
  signal tmp_ivl_39607 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4783
  signal tmp_ivl_39609 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4783
  signal tmp_ivl_39614 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4783
  signal tmp_ivl_39617 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4783
  signal tmp_ivl_39621 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4783
  signal tmp_ivl_39623 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4783
  signal tmp_ivl_39625 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4783
  signal tmp_ivl_39631 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4784
  signal tmp_ivl_39632 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4784
  signal tmp_ivl_39637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4784
  signal tmp_ivl_39639 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4784
  signal tmp_ivl_3964 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3077
  signal tmp_ivl_39644 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4784
  signal tmp_ivl_39647 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4784
  signal tmp_ivl_39651 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4784
  signal tmp_ivl_39653 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4784
  signal tmp_ivl_39655 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4784
  signal tmp_ivl_39661 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4785
  signal tmp_ivl_39662 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4785
  signal tmp_ivl_39667 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4785
  signal tmp_ivl_39669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4785
  signal tmp_ivl_3967 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3077
  signal tmp_ivl_39674 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4785
  signal tmp_ivl_39677 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4785
  signal tmp_ivl_39681 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4785
  signal tmp_ivl_39683 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4785
  signal tmp_ivl_39685 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4785
  signal tmp_ivl_3969 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3077
  signal tmp_ivl_39691 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4786
  signal tmp_ivl_39692 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4786
  signal tmp_ivl_39697 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4786
  signal tmp_ivl_39699 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4786
  signal tmp_ivl_397 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2953
  signal tmp_ivl_3970 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3077
  signal tmp_ivl_39704 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4786
  signal tmp_ivl_39707 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4786
  signal tmp_ivl_39711 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4786
  signal tmp_ivl_39713 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4786
  signal tmp_ivl_39715 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4786
  signal tmp_ivl_39721 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4787
  signal tmp_ivl_39722 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4787
  signal tmp_ivl_39727 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4787
  signal tmp_ivl_39729 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4787
  signal tmp_ivl_39734 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4787
  signal tmp_ivl_39737 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4787
  signal tmp_ivl_39741 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4787
  signal tmp_ivl_39743 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4787
  signal tmp_ivl_39745 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4787
  signal tmp_ivl_3975 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3077
  signal tmp_ivl_39751 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4788
  signal tmp_ivl_39752 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4788
  signal tmp_ivl_39757 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4788
  signal tmp_ivl_39759 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4788
  signal tmp_ivl_39764 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4788
  signal tmp_ivl_39767 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4788
  signal tmp_ivl_3977 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3077
  signal tmp_ivl_39771 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4788
  signal tmp_ivl_39773 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4788
  signal tmp_ivl_39775 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4788
  signal tmp_ivl_39781 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4789
  signal tmp_ivl_39782 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4789
  signal tmp_ivl_39787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4789
  signal tmp_ivl_39789 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4789
  signal tmp_ivl_39794 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4789
  signal tmp_ivl_39797 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4789
  signal tmp_ivl_39801 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4789
  signal tmp_ivl_39803 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4789
  signal tmp_ivl_39805 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4789
  signal tmp_ivl_39811 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4790
  signal tmp_ivl_39812 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4790
  signal tmp_ivl_39817 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4790
  signal tmp_ivl_39819 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4790
  signal tmp_ivl_39824 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4790
  signal tmp_ivl_39827 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4790
  signal tmp_ivl_3983 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3078
  signal tmp_ivl_39831 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4790
  signal tmp_ivl_39833 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4790
  signal tmp_ivl_39835 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4790
  signal tmp_ivl_39841 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4791
  signal tmp_ivl_39842 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4791
  signal tmp_ivl_39847 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4791
  signal tmp_ivl_39849 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4791
  signal tmp_ivl_3985 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3078
  signal tmp_ivl_39854 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4791
  signal tmp_ivl_39857 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4791
  signal tmp_ivl_3986 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3078
  signal tmp_ivl_39861 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4791
  signal tmp_ivl_39863 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4791
  signal tmp_ivl_39865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4791
  signal tmp_ivl_39871 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4792
  signal tmp_ivl_39872 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4792
  signal tmp_ivl_39877 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4792
  signal tmp_ivl_39879 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4792
  signal tmp_ivl_39884 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4792
  signal tmp_ivl_39887 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4792
  signal tmp_ivl_39891 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4792
  signal tmp_ivl_39893 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4792
  signal tmp_ivl_39895 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4792
  signal tmp_ivl_399 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2953
  signal tmp_ivl_39901 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4793
  signal tmp_ivl_39902 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4793
  signal tmp_ivl_39907 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4793
  signal tmp_ivl_39909 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4793
  signal tmp_ivl_3991 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3078
  signal tmp_ivl_39914 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4793
  signal tmp_ivl_39917 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4793
  signal tmp_ivl_39921 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4793
  signal tmp_ivl_39923 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4793
  signal tmp_ivl_39925 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4793
  signal tmp_ivl_39931 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4794
  signal tmp_ivl_39932 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4794
  signal tmp_ivl_39937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4794
  signal tmp_ivl_39939 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4794
  signal tmp_ivl_3994 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3078
  signal tmp_ivl_39944 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4794
  signal tmp_ivl_39947 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4794
  signal tmp_ivl_39951 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4794
  signal tmp_ivl_39953 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4794
  signal tmp_ivl_39955 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4794
  signal tmp_ivl_3996 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3078
  signal tmp_ivl_39961 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4795
  signal tmp_ivl_39962 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4795
  signal tmp_ivl_39967 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4795
  signal tmp_ivl_39969 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4795
  signal tmp_ivl_3997 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3078
  signal tmp_ivl_39974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4795
  signal tmp_ivl_39977 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4795
  signal tmp_ivl_39981 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4795
  signal tmp_ivl_39983 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4795
  signal tmp_ivl_39985 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4795
  signal tmp_ivl_39991 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4796
  signal tmp_ivl_39992 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4796
  signal tmp_ivl_39997 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4796
  signal tmp_ivl_39999 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4796
  signal tmp_ivl_4 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2940
  signal tmp_ivl_40004 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4796
  signal tmp_ivl_40007 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4796
  signal tmp_ivl_40011 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4796
  signal tmp_ivl_40013 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4796
  signal tmp_ivl_40015 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4796
  signal tmp_ivl_4002 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3078
  signal tmp_ivl_40021 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4797
  signal tmp_ivl_40022 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4797
  signal tmp_ivl_40027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4797
  signal tmp_ivl_40029 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4797
  signal tmp_ivl_40034 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4797
  signal tmp_ivl_40037 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4797
  signal tmp_ivl_4004 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3078
  signal tmp_ivl_40041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4797
  signal tmp_ivl_40043 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4797
  signal tmp_ivl_40045 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4797
  signal tmp_ivl_40051 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4798
  signal tmp_ivl_40052 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4798
  signal tmp_ivl_40057 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4798
  signal tmp_ivl_40059 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4798
  signal tmp_ivl_40064 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4798
  signal tmp_ivl_40067 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4798
  signal tmp_ivl_40071 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4798
  signal tmp_ivl_40073 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4798
  signal tmp_ivl_40075 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4798
  signal tmp_ivl_40081 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4799
  signal tmp_ivl_40082 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4799
  signal tmp_ivl_40087 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4799
  signal tmp_ivl_40089 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4799
  signal tmp_ivl_40094 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4799
  signal tmp_ivl_40097 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4799
  signal tmp_ivl_401 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2953
  signal tmp_ivl_4010 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3079
  signal tmp_ivl_40101 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4799
  signal tmp_ivl_40103 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4799
  signal tmp_ivl_40105 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4799
  signal tmp_ivl_40111 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4800
  signal tmp_ivl_40112 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4800
  signal tmp_ivl_40117 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4800
  signal tmp_ivl_40119 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4800
  signal tmp_ivl_4012 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3079
  signal tmp_ivl_40124 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4800
  signal tmp_ivl_40127 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4800
  signal tmp_ivl_4013 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3079
  signal tmp_ivl_40131 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4800
  signal tmp_ivl_40133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4800
  signal tmp_ivl_40135 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4800
  signal tmp_ivl_40141 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4801
  signal tmp_ivl_40142 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4801
  signal tmp_ivl_40147 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4801
  signal tmp_ivl_40149 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4801
  signal tmp_ivl_40154 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4801
  signal tmp_ivl_40157 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4801
  signal tmp_ivl_40161 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4801
  signal tmp_ivl_40163 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4801
  signal tmp_ivl_40165 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4801
  signal tmp_ivl_40171 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4802
  signal tmp_ivl_40172 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4802
  signal tmp_ivl_40177 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4802
  signal tmp_ivl_40179 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4802
  signal tmp_ivl_4018 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3079
  signal tmp_ivl_40184 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4802
  signal tmp_ivl_40187 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4802
  signal tmp_ivl_40191 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4802
  signal tmp_ivl_40193 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4802
  signal tmp_ivl_40195 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4802
  signal tmp_ivl_40201 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4803
  signal tmp_ivl_40202 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4803
  signal tmp_ivl_40207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4803
  signal tmp_ivl_40209 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4803
  signal tmp_ivl_4021 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3079
  signal tmp_ivl_40214 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4803
  signal tmp_ivl_40217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4803
  signal tmp_ivl_40221 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4803
  signal tmp_ivl_40223 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4803
  signal tmp_ivl_40225 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4803
  signal tmp_ivl_4023 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3079
  signal tmp_ivl_40231 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4804
  signal tmp_ivl_40232 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4804
  signal tmp_ivl_40237 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4804
  signal tmp_ivl_40239 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4804
  signal tmp_ivl_4024 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3079
  signal tmp_ivl_40244 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4804
  signal tmp_ivl_40247 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4804
  signal tmp_ivl_40251 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4804
  signal tmp_ivl_40253 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4804
  signal tmp_ivl_40255 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4804
  signal tmp_ivl_40261 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4805
  signal tmp_ivl_40262 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4805
  signal tmp_ivl_40267 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4805
  signal tmp_ivl_40269 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4805
  signal tmp_ivl_40274 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4805
  signal tmp_ivl_40277 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4805
  signal tmp_ivl_40281 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4805
  signal tmp_ivl_40283 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4805
  signal tmp_ivl_40285 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4805
  signal tmp_ivl_4029 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3079
  signal tmp_ivl_40291 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4806
  signal tmp_ivl_40292 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4806
  signal tmp_ivl_40297 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4806
  signal tmp_ivl_40299 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4806
  signal tmp_ivl_40304 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4806
  signal tmp_ivl_40307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4806
  signal tmp_ivl_4031 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3079
  signal tmp_ivl_40311 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4806
  signal tmp_ivl_40313 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4806
  signal tmp_ivl_40315 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4806
  signal tmp_ivl_40321 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4807
  signal tmp_ivl_40322 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4807
  signal tmp_ivl_40327 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4807
  signal tmp_ivl_40329 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4807
  signal tmp_ivl_40334 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4807
  signal tmp_ivl_40337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4807
  signal tmp_ivl_40341 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4807
  signal tmp_ivl_40343 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4807
  signal tmp_ivl_40345 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4807
  signal tmp_ivl_40351 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4808
  signal tmp_ivl_40352 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4808
  signal tmp_ivl_40357 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4808
  signal tmp_ivl_40359 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4808
  signal tmp_ivl_40364 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4808
  signal tmp_ivl_40367 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4808
  signal tmp_ivl_4037 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3080
  signal tmp_ivl_40371 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4808
  signal tmp_ivl_40373 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4808
  signal tmp_ivl_40375 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4808
  signal tmp_ivl_40381 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4809
  signal tmp_ivl_40382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4809
  signal tmp_ivl_40387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4809
  signal tmp_ivl_40389 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4809
  signal tmp_ivl_4039 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3080
  signal tmp_ivl_40394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4809
  signal tmp_ivl_40397 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4809
  signal tmp_ivl_4040 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3080
  signal tmp_ivl_40401 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4809
  signal tmp_ivl_40403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4809
  signal tmp_ivl_40405 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4809
  signal tmp_ivl_40411 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4810
  signal tmp_ivl_40412 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4810
  signal tmp_ivl_40417 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4810
  signal tmp_ivl_40419 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4810
  signal tmp_ivl_40424 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4810
  signal tmp_ivl_40427 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4810
  signal tmp_ivl_40431 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4810
  signal tmp_ivl_40433 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4810
  signal tmp_ivl_40435 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4810
  signal tmp_ivl_40441 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4811
  signal tmp_ivl_40442 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4811
  signal tmp_ivl_40447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4811
  signal tmp_ivl_40449 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4811
  signal tmp_ivl_4045 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3080
  signal tmp_ivl_40454 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4811
  signal tmp_ivl_40457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4811
  signal tmp_ivl_40461 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4811
  signal tmp_ivl_40463 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4811
  signal tmp_ivl_40465 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4811
  signal tmp_ivl_40471 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4812
  signal tmp_ivl_40472 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4812
  signal tmp_ivl_40477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4812
  signal tmp_ivl_40479 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4812
  signal tmp_ivl_4048 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3080
  signal tmp_ivl_40484 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4812
  signal tmp_ivl_40487 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4812
  signal tmp_ivl_40491 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4812
  signal tmp_ivl_40493 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4812
  signal tmp_ivl_40495 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4812
  signal tmp_ivl_4050 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3080
  signal tmp_ivl_40501 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4813
  signal tmp_ivl_40502 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4813
  signal tmp_ivl_40507 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4813
  signal tmp_ivl_40509 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4813
  signal tmp_ivl_4051 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3080
  signal tmp_ivl_40514 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4813
  signal tmp_ivl_40517 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4813
  signal tmp_ivl_40521 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4813
  signal tmp_ivl_40523 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4813
  signal tmp_ivl_40525 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4813
  signal tmp_ivl_40531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4814
  signal tmp_ivl_40532 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4814
  signal tmp_ivl_40537 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4814
  signal tmp_ivl_40539 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4814
  signal tmp_ivl_40544 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4814
  signal tmp_ivl_40547 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4814
  signal tmp_ivl_40551 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4814
  signal tmp_ivl_40553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4814
  signal tmp_ivl_40555 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4814
  signal tmp_ivl_4056 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3080
  signal tmp_ivl_40561 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4815
  signal tmp_ivl_40562 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4815
  signal tmp_ivl_40567 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4815
  signal tmp_ivl_40569 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4815
  signal tmp_ivl_40574 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4815
  signal tmp_ivl_40577 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4815
  signal tmp_ivl_4058 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3080
  signal tmp_ivl_40581 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4815
  signal tmp_ivl_40583 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4815
  signal tmp_ivl_40585 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4815
  signal tmp_ivl_40591 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4816
  signal tmp_ivl_40592 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4816
  signal tmp_ivl_40597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4816
  signal tmp_ivl_40599 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4816
  signal tmp_ivl_40604 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4816
  signal tmp_ivl_40607 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4816
  signal tmp_ivl_40611 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4816
  signal tmp_ivl_40613 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4816
  signal tmp_ivl_40615 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4816
  signal tmp_ivl_40621 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4817
  signal tmp_ivl_40622 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4817
  signal tmp_ivl_40627 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4817
  signal tmp_ivl_40629 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4817
  signal tmp_ivl_40634 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4817
  signal tmp_ivl_40637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4817
  signal tmp_ivl_4064 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3081
  signal tmp_ivl_40641 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4817
  signal tmp_ivl_40643 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4817
  signal tmp_ivl_40645 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4817
  signal tmp_ivl_40651 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4818
  signal tmp_ivl_40652 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4818
  signal tmp_ivl_40657 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4818
  signal tmp_ivl_40659 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4818
  signal tmp_ivl_4066 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3081
  signal tmp_ivl_40664 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4818
  signal tmp_ivl_40667 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4818
  signal tmp_ivl_4067 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3081
  signal tmp_ivl_40671 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4818
  signal tmp_ivl_40673 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4818
  signal tmp_ivl_40675 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4818
  signal tmp_ivl_40681 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4819
  signal tmp_ivl_40682 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4819
  signal tmp_ivl_40687 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4819
  signal tmp_ivl_40689 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4819
  signal tmp_ivl_40694 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4819
  signal tmp_ivl_40697 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4819
  signal tmp_ivl_407 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2954
  signal tmp_ivl_40701 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4819
  signal tmp_ivl_40703 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4819
  signal tmp_ivl_40705 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4819
  signal tmp_ivl_40711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4820
  signal tmp_ivl_40712 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4820
  signal tmp_ivl_40717 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4820
  signal tmp_ivl_40719 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4820
  signal tmp_ivl_4072 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3081
  signal tmp_ivl_40724 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4820
  signal tmp_ivl_40727 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4820
  signal tmp_ivl_40731 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4820
  signal tmp_ivl_40733 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4820
  signal tmp_ivl_40735 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4820
  signal tmp_ivl_40741 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4821
  signal tmp_ivl_40742 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4821
  signal tmp_ivl_40747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4821
  signal tmp_ivl_40749 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4821
  signal tmp_ivl_4075 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3081
  signal tmp_ivl_40754 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4821
  signal tmp_ivl_40757 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4821
  signal tmp_ivl_40761 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4821
  signal tmp_ivl_40763 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4821
  signal tmp_ivl_40765 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4821
  signal tmp_ivl_4077 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3081
  signal tmp_ivl_40770 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4822
  signal tmp_ivl_40775 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4822
  signal tmp_ivl_40778 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4822
  signal tmp_ivl_40779 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4822
  signal tmp_ivl_4078 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3081
  signal tmp_ivl_40784 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4822
  signal tmp_ivl_40787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4822
  signal tmp_ivl_40791 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4822
  signal tmp_ivl_40793 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4822
  signal tmp_ivl_40795 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4822
  signal tmp_ivl_40800 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4823
  signal tmp_ivl_40805 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4823
  signal tmp_ivl_40808 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4823
  signal tmp_ivl_40809 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4823
  signal tmp_ivl_40814 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4823
  signal tmp_ivl_40817 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4823
  signal tmp_ivl_40821 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4823
  signal tmp_ivl_40823 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4823
  signal tmp_ivl_40825 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4823
  signal tmp_ivl_4083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3081
  signal tmp_ivl_40830 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4824
  signal tmp_ivl_40835 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4824
  signal tmp_ivl_40838 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4824
  signal tmp_ivl_40839 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4824
  signal tmp_ivl_40844 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4824
  signal tmp_ivl_40847 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4824
  signal tmp_ivl_4085 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3081
  signal tmp_ivl_40851 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4824
  signal tmp_ivl_40853 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4824
  signal tmp_ivl_40855 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4824
  signal tmp_ivl_40860 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4825
  signal tmp_ivl_40865 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4825
  signal tmp_ivl_40868 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4825
  signal tmp_ivl_40869 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4825
  signal tmp_ivl_40874 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4825
  signal tmp_ivl_40877 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4825
  signal tmp_ivl_40881 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4825
  signal tmp_ivl_40883 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4825
  signal tmp_ivl_40885 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4825
  signal tmp_ivl_40890 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4826
  signal tmp_ivl_40895 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4826
  signal tmp_ivl_40898 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4826
  signal tmp_ivl_40899 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4826
  signal tmp_ivl_409 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2954
  signal tmp_ivl_40904 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4826
  signal tmp_ivl_40907 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4826
  signal tmp_ivl_4091 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3082
  signal tmp_ivl_40911 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4826
  signal tmp_ivl_40913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4826
  signal tmp_ivl_40915 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4826
  signal tmp_ivl_40920 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4827
  signal tmp_ivl_40925 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4827
  signal tmp_ivl_40928 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4827
  signal tmp_ivl_40929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4827
  signal tmp_ivl_4093 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3082
  signal tmp_ivl_40934 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4827
  signal tmp_ivl_40937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4827
  signal tmp_ivl_4094 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3082
  signal tmp_ivl_40941 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4827
  signal tmp_ivl_40943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4827
  signal tmp_ivl_40945 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4827
  signal tmp_ivl_40950 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4828
  signal tmp_ivl_40955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4828
  signal tmp_ivl_40958 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4828
  signal tmp_ivl_40959 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4828
  signal tmp_ivl_40964 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4828
  signal tmp_ivl_40967 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4828
  signal tmp_ivl_40971 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4828
  signal tmp_ivl_40973 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4828
  signal tmp_ivl_40975 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4828
  signal tmp_ivl_40980 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4829
  signal tmp_ivl_40985 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4829
  signal tmp_ivl_40988 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4829
  signal tmp_ivl_40989 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4829
  signal tmp_ivl_4099 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3082
  signal tmp_ivl_40994 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4829
  signal tmp_ivl_40997 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4829
  signal tmp_ivl_41 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2941
  signal tmp_ivl_410 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2954
  signal tmp_ivl_41001 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4829
  signal tmp_ivl_41003 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4829
  signal tmp_ivl_41005 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4829
  signal tmp_ivl_41010 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4830
  signal tmp_ivl_41015 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4830
  signal tmp_ivl_41018 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4830
  signal tmp_ivl_41019 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4830
  signal tmp_ivl_4102 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3082
  signal tmp_ivl_41024 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4830
  signal tmp_ivl_41027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4830
  signal tmp_ivl_41031 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4830
  signal tmp_ivl_41033 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4830
  signal tmp_ivl_41035 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4830
  signal tmp_ivl_4104 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3082
  signal tmp_ivl_41040 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4831
  signal tmp_ivl_41045 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4831
  signal tmp_ivl_41048 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4831
  signal tmp_ivl_41049 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4831
  signal tmp_ivl_4105 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3082
  signal tmp_ivl_41054 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4831
  signal tmp_ivl_41057 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4831
  signal tmp_ivl_41061 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4831
  signal tmp_ivl_41063 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4831
  signal tmp_ivl_41065 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4831
  signal tmp_ivl_41070 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4832
  signal tmp_ivl_41075 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4832
  signal tmp_ivl_41078 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4832
  signal tmp_ivl_41079 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4832
  signal tmp_ivl_41084 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4832
  signal tmp_ivl_41087 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4832
  signal tmp_ivl_41091 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4832
  signal tmp_ivl_41093 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4832
  signal tmp_ivl_41095 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4832
  signal tmp_ivl_4110 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3082
  signal tmp_ivl_41100 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4833
  signal tmp_ivl_41105 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4833
  signal tmp_ivl_41108 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4833
  signal tmp_ivl_41109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4833
  signal tmp_ivl_41114 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4833
  signal tmp_ivl_41117 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4833
  signal tmp_ivl_4112 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3082
  signal tmp_ivl_41121 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4833
  signal tmp_ivl_41123 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4833
  signal tmp_ivl_41125 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4833
  signal tmp_ivl_41130 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4834
  signal tmp_ivl_41135 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4834
  signal tmp_ivl_41138 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4834
  signal tmp_ivl_41139 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4834
  signal tmp_ivl_41144 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4834
  signal tmp_ivl_41147 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4834
  signal tmp_ivl_41151 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4834
  signal tmp_ivl_41153 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4834
  signal tmp_ivl_41155 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4834
  signal tmp_ivl_41160 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4835
  signal tmp_ivl_41165 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4835
  signal tmp_ivl_41168 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4835
  signal tmp_ivl_41169 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4835
  signal tmp_ivl_41174 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4835
  signal tmp_ivl_41177 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4835
  signal tmp_ivl_4118 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3083
  signal tmp_ivl_41181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4835
  signal tmp_ivl_41183 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4835
  signal tmp_ivl_41185 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4835
  signal tmp_ivl_41190 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4836
  signal tmp_ivl_41195 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4836
  signal tmp_ivl_41198 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4836
  signal tmp_ivl_41199 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4836
  signal tmp_ivl_4120 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3083
  signal tmp_ivl_41204 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4836
  signal tmp_ivl_41207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4836
  signal tmp_ivl_4121 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3083
  signal tmp_ivl_41211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4836
  signal tmp_ivl_41213 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4836
  signal tmp_ivl_41215 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4836
  signal tmp_ivl_41220 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4837
  signal tmp_ivl_41225 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4837
  signal tmp_ivl_41228 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4837
  signal tmp_ivl_41229 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4837
  signal tmp_ivl_41234 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4837
  signal tmp_ivl_41237 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4837
  signal tmp_ivl_41241 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4837
  signal tmp_ivl_41243 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4837
  signal tmp_ivl_41245 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4837
  signal tmp_ivl_41250 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4838
  signal tmp_ivl_41255 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4838
  signal tmp_ivl_41258 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4838
  signal tmp_ivl_41259 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4838
  signal tmp_ivl_4126 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3083
  signal tmp_ivl_41264 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4838
  signal tmp_ivl_41267 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4838
  signal tmp_ivl_41271 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4838
  signal tmp_ivl_41273 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4838
  signal tmp_ivl_41275 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4838
  signal tmp_ivl_41280 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4839
  signal tmp_ivl_41285 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4839
  signal tmp_ivl_41288 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4839
  signal tmp_ivl_41289 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4839
  signal tmp_ivl_4129 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3083
  signal tmp_ivl_41294 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4839
  signal tmp_ivl_41297 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4839
  signal tmp_ivl_41301 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4839
  signal tmp_ivl_41303 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4839
  signal tmp_ivl_41305 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4839
  signal tmp_ivl_4131 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3083
  signal tmp_ivl_41310 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4840
  signal tmp_ivl_41315 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4840
  signal tmp_ivl_41318 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4840
  signal tmp_ivl_41319 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4840
  signal tmp_ivl_4132 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3083
  signal tmp_ivl_41324 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4840
  signal tmp_ivl_41327 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4840
  signal tmp_ivl_41331 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4840
  signal tmp_ivl_41333 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4840
  signal tmp_ivl_41335 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4840
  signal tmp_ivl_41340 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4841
  signal tmp_ivl_41345 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4841
  signal tmp_ivl_41348 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4841
  signal tmp_ivl_41349 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4841
  signal tmp_ivl_41354 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4841
  signal tmp_ivl_41357 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4841
  signal tmp_ivl_41361 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4841
  signal tmp_ivl_41363 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4841
  signal tmp_ivl_41365 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4841
  signal tmp_ivl_4137 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3083
  signal tmp_ivl_41370 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4842
  signal tmp_ivl_41375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4842
  signal tmp_ivl_41378 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4842
  signal tmp_ivl_41379 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4842
  signal tmp_ivl_41384 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4842
  signal tmp_ivl_41387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4842
  signal tmp_ivl_4139 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3083
  signal tmp_ivl_41391 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4842
  signal tmp_ivl_41393 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4842
  signal tmp_ivl_41395 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4842
  signal tmp_ivl_41400 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4843
  signal tmp_ivl_41405 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4843
  signal tmp_ivl_41408 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4843
  signal tmp_ivl_41409 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4843
  signal tmp_ivl_41414 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4843
  signal tmp_ivl_41417 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4843
  signal tmp_ivl_41421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4843
  signal tmp_ivl_41423 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4843
  signal tmp_ivl_41425 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4843
  signal tmp_ivl_41430 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4844
  signal tmp_ivl_41435 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4844
  signal tmp_ivl_41438 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4844
  signal tmp_ivl_41439 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4844
  signal tmp_ivl_41444 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4844
  signal tmp_ivl_41447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4844
  signal tmp_ivl_4145 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3084
  signal tmp_ivl_41451 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4844
  signal tmp_ivl_41453 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4844
  signal tmp_ivl_41455 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4844
  signal tmp_ivl_41460 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4845
  signal tmp_ivl_41465 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4845
  signal tmp_ivl_41468 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4845
  signal tmp_ivl_41469 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4845
  signal tmp_ivl_4147 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3084
  signal tmp_ivl_41474 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4845
  signal tmp_ivl_41477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4845
  signal tmp_ivl_4148 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3084
  signal tmp_ivl_41481 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4845
  signal tmp_ivl_41483 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4845
  signal tmp_ivl_41485 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4845
  signal tmp_ivl_41490 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4846
  signal tmp_ivl_41495 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4846
  signal tmp_ivl_41498 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4846
  signal tmp_ivl_41499 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4846
  signal tmp_ivl_415 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2954
  signal tmp_ivl_41504 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4846
  signal tmp_ivl_41507 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4846
  signal tmp_ivl_41511 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4846
  signal tmp_ivl_41513 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4846
  signal tmp_ivl_41515 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4846
  signal tmp_ivl_41520 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4847
  signal tmp_ivl_41525 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4847
  signal tmp_ivl_41528 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4847
  signal tmp_ivl_41529 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4847
  signal tmp_ivl_4153 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3084
  signal tmp_ivl_41534 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4847
  signal tmp_ivl_41537 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4847
  signal tmp_ivl_41541 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4847
  signal tmp_ivl_41543 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4847
  signal tmp_ivl_41545 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4847
  signal tmp_ivl_41550 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4848
  signal tmp_ivl_41555 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4848
  signal tmp_ivl_41558 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4848
  signal tmp_ivl_41559 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4848
  signal tmp_ivl_4156 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3084
  signal tmp_ivl_41564 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4848
  signal tmp_ivl_41567 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4848
  signal tmp_ivl_41571 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4848
  signal tmp_ivl_41573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4848
  signal tmp_ivl_41575 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4848
  signal tmp_ivl_4158 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3084
  signal tmp_ivl_41580 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4849
  signal tmp_ivl_41585 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4849
  signal tmp_ivl_41588 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4849
  signal tmp_ivl_41589 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4849
  signal tmp_ivl_4159 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3084
  signal tmp_ivl_41594 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4849
  signal tmp_ivl_41597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4849
  signal tmp_ivl_41601 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4849
  signal tmp_ivl_41603 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4849
  signal tmp_ivl_41605 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4849
  signal tmp_ivl_41610 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4850
  signal tmp_ivl_41615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4850
  signal tmp_ivl_41618 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4850
  signal tmp_ivl_41619 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4850
  signal tmp_ivl_41624 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4850
  signal tmp_ivl_41627 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4850
  signal tmp_ivl_41631 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4850
  signal tmp_ivl_41633 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4850
  signal tmp_ivl_41635 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4850
  signal tmp_ivl_4164 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3084
  signal tmp_ivl_41640 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4851
  signal tmp_ivl_41645 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4851
  signal tmp_ivl_41648 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4851
  signal tmp_ivl_41649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4851
  signal tmp_ivl_41654 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4851
  signal tmp_ivl_41657 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4851
  signal tmp_ivl_4166 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3084
  signal tmp_ivl_41661 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4851
  signal tmp_ivl_41663 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4851
  signal tmp_ivl_41665 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4851
  signal tmp_ivl_41670 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4852
  signal tmp_ivl_41675 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4852
  signal tmp_ivl_41678 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4852
  signal tmp_ivl_41679 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4852
  signal tmp_ivl_41684 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4852
  signal tmp_ivl_41687 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4852
  signal tmp_ivl_41691 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4852
  signal tmp_ivl_41693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4852
  signal tmp_ivl_41695 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4852
  signal tmp_ivl_41700 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4853
  signal tmp_ivl_41705 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4853
  signal tmp_ivl_41708 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4853
  signal tmp_ivl_41709 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4853
  signal tmp_ivl_41714 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4853
  signal tmp_ivl_41717 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4853
  signal tmp_ivl_4172 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3085
  signal tmp_ivl_41721 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4853
  signal tmp_ivl_41723 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4853
  signal tmp_ivl_41725 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4853
  signal tmp_ivl_41730 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4854
  signal tmp_ivl_41735 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4854
  signal tmp_ivl_41738 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4854
  signal tmp_ivl_41739 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4854
  signal tmp_ivl_4174 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3085
  signal tmp_ivl_41744 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4854
  signal tmp_ivl_41747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4854
  signal tmp_ivl_4175 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3085
  signal tmp_ivl_41751 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4854
  signal tmp_ivl_41753 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4854
  signal tmp_ivl_41755 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4854
  signal tmp_ivl_41760 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4855
  signal tmp_ivl_41765 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4855
  signal tmp_ivl_41768 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4855
  signal tmp_ivl_41769 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4855
  signal tmp_ivl_41774 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4855
  signal tmp_ivl_41777 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4855
  signal tmp_ivl_41781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4855
  signal tmp_ivl_41783 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4855
  signal tmp_ivl_41785 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4855
  signal tmp_ivl_41790 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4856
  signal tmp_ivl_41795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4856
  signal tmp_ivl_41798 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4856
  signal tmp_ivl_41799 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4856
  signal tmp_ivl_418 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2954
  signal tmp_ivl_4180 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3085
  signal tmp_ivl_41804 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4856
  signal tmp_ivl_41807 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4856
  signal tmp_ivl_41811 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4856
  signal tmp_ivl_41813 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4856
  signal tmp_ivl_41815 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4856
  signal tmp_ivl_41820 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4857
  signal tmp_ivl_41825 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4857
  signal tmp_ivl_41828 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4857
  signal tmp_ivl_41829 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4857
  signal tmp_ivl_4183 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3085
  signal tmp_ivl_41834 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4857
  signal tmp_ivl_41837 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4857
  signal tmp_ivl_41841 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4857
  signal tmp_ivl_41843 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4857
  signal tmp_ivl_41845 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4857
  signal tmp_ivl_4185 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3085
  signal tmp_ivl_41850 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4858
  signal tmp_ivl_41855 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4858
  signal tmp_ivl_41858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4858
  signal tmp_ivl_41859 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4858
  signal tmp_ivl_4186 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3085
  signal tmp_ivl_41864 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4858
  signal tmp_ivl_41867 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4858
  signal tmp_ivl_41871 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4858
  signal tmp_ivl_41873 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4858
  signal tmp_ivl_41875 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4858
  signal tmp_ivl_41880 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4859
  signal tmp_ivl_41885 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4859
  signal tmp_ivl_41888 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4859
  signal tmp_ivl_41889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4859
  signal tmp_ivl_41894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4859
  signal tmp_ivl_41897 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4859
  signal tmp_ivl_41901 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4859
  signal tmp_ivl_41903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4859
  signal tmp_ivl_41905 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4859
  signal tmp_ivl_4191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3085
  signal tmp_ivl_41910 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4860
  signal tmp_ivl_41915 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4860
  signal tmp_ivl_41917 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4860
  signal tmp_ivl_41922 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4860
  signal tmp_ivl_41925 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4860
  signal tmp_ivl_41929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4860
  signal tmp_ivl_4193 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3085
  signal tmp_ivl_41931 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4860
  signal tmp_ivl_41933 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4860
  signal tmp_ivl_41938 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4861
  signal tmp_ivl_41943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4861
  signal tmp_ivl_41945 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4861
  signal tmp_ivl_41950 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4861
  signal tmp_ivl_41953 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4861
  signal tmp_ivl_41957 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4861
  signal tmp_ivl_41959 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4861
  signal tmp_ivl_41961 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4861
  signal tmp_ivl_41966 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4862
  signal tmp_ivl_41971 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4862
  signal tmp_ivl_41973 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4862
  signal tmp_ivl_41978 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4862
  signal tmp_ivl_41981 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4862
  signal tmp_ivl_41985 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4862
  signal tmp_ivl_41987 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4862
  signal tmp_ivl_41989 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4862
  signal tmp_ivl_4199 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3086
  signal tmp_ivl_41994 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4863
  signal tmp_ivl_41999 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4863
  signal tmp_ivl_420 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2954
  signal tmp_ivl_42001 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4863
  signal tmp_ivl_42006 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4863
  signal tmp_ivl_42009 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4863
  signal tmp_ivl_4201 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3086
  signal tmp_ivl_42013 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4863
  signal tmp_ivl_42015 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4863
  signal tmp_ivl_42017 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4863
  signal tmp_ivl_4202 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3086
  signal tmp_ivl_42022 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4864
  signal tmp_ivl_42027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4864
  signal tmp_ivl_42029 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4864
  signal tmp_ivl_42034 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4864
  signal tmp_ivl_42037 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4864
  signal tmp_ivl_42041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4864
  signal tmp_ivl_42043 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4864
  signal tmp_ivl_42045 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4864
  signal tmp_ivl_42050 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4865
  signal tmp_ivl_42055 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4865
  signal tmp_ivl_42057 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4865
  signal tmp_ivl_42062 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4865
  signal tmp_ivl_42065 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4865
  signal tmp_ivl_42069 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4865
  signal tmp_ivl_4207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3086
  signal tmp_ivl_42071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4865
  signal tmp_ivl_42073 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4865
  signal tmp_ivl_42078 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4866
  signal tmp_ivl_42083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4866
  signal tmp_ivl_42085 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4866
  signal tmp_ivl_42090 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4866
  signal tmp_ivl_42093 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4866
  signal tmp_ivl_42097 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4866
  signal tmp_ivl_42099 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4866
  signal tmp_ivl_421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2954
  signal tmp_ivl_4210 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3086
  signal tmp_ivl_42101 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4866
  signal tmp_ivl_42106 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4867
  signal tmp_ivl_42111 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4867
  signal tmp_ivl_42113 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4867
  signal tmp_ivl_42118 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4867
  signal tmp_ivl_4212 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3086
  signal tmp_ivl_42121 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4867
  signal tmp_ivl_42125 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4867
  signal tmp_ivl_42127 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4867
  signal tmp_ivl_42129 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4867
  signal tmp_ivl_4213 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3086
  signal tmp_ivl_42134 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4868
  signal tmp_ivl_42139 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4868
  signal tmp_ivl_42141 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4868
  signal tmp_ivl_42146 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4868
  signal tmp_ivl_42149 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4868
  signal tmp_ivl_42153 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4868
  signal tmp_ivl_42155 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4868
  signal tmp_ivl_42157 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4868
  signal tmp_ivl_42162 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4869
  signal tmp_ivl_42167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4869
  signal tmp_ivl_42169 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4869
  signal tmp_ivl_42174 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4869
  signal tmp_ivl_42177 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4869
  signal tmp_ivl_4218 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3086
  signal tmp_ivl_42181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4869
  signal tmp_ivl_42183 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4869
  signal tmp_ivl_42185 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4869
  signal tmp_ivl_42191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4870
  signal tmp_ivl_42192 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4870
  signal tmp_ivl_42197 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4870
  signal tmp_ivl_42199 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4870
  signal tmp_ivl_4220 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3086
  signal tmp_ivl_42204 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4870
  signal tmp_ivl_42207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4870
  signal tmp_ivl_42211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4870
  signal tmp_ivl_42213 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4870
  signal tmp_ivl_42215 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4870
  signal tmp_ivl_42220 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4871
  signal tmp_ivl_42225 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4871
  signal tmp_ivl_42227 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4871
  signal tmp_ivl_42232 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4871
  signal tmp_ivl_42235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4871
  signal tmp_ivl_42239 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4871
  signal tmp_ivl_42241 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4871
  signal tmp_ivl_42243 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4871
  signal tmp_ivl_42249 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4872
  signal tmp_ivl_42250 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4872
  signal tmp_ivl_42255 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4872
  signal tmp_ivl_42257 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4872
  signal tmp_ivl_4226 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3087
  signal tmp_ivl_42262 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4872
  signal tmp_ivl_42265 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4872
  signal tmp_ivl_42269 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4872
  signal tmp_ivl_42271 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4872
  signal tmp_ivl_42273 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4872
  signal tmp_ivl_42278 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4873
  signal tmp_ivl_4228 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3087
  signal tmp_ivl_42283 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4873
  signal tmp_ivl_42285 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4873
  signal tmp_ivl_4229 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3087
  signal tmp_ivl_42290 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4873
  signal tmp_ivl_42293 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4873
  signal tmp_ivl_42297 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4873
  signal tmp_ivl_42299 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4873
  signal tmp_ivl_42301 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4873
  signal tmp_ivl_42306 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4874
  signal tmp_ivl_42311 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4874
  signal tmp_ivl_42313 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4874
  signal tmp_ivl_42318 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4874
  signal tmp_ivl_42321 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4874
  signal tmp_ivl_42325 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4874
  signal tmp_ivl_42327 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4874
  signal tmp_ivl_42329 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4874
  signal tmp_ivl_42334 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4875
  signal tmp_ivl_42339 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4875
  signal tmp_ivl_4234 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3087
  signal tmp_ivl_42341 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4875
  signal tmp_ivl_42346 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4875
  signal tmp_ivl_42349 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4875
  signal tmp_ivl_42353 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4875
  signal tmp_ivl_42355 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4875
  signal tmp_ivl_42357 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4875
  signal tmp_ivl_42362 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4876
  signal tmp_ivl_42367 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4876
  signal tmp_ivl_42369 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4876
  signal tmp_ivl_4237 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3087
  signal tmp_ivl_42374 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4876
  signal tmp_ivl_42377 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4876
  signal tmp_ivl_42381 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4876
  signal tmp_ivl_42383 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4876
  signal tmp_ivl_42385 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4876
  signal tmp_ivl_4239 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3087
  signal tmp_ivl_42390 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4877
  signal tmp_ivl_42395 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4877
  signal tmp_ivl_42397 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4877
  signal tmp_ivl_4240 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3087
  signal tmp_ivl_42402 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4877
  signal tmp_ivl_42405 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4877
  signal tmp_ivl_42409 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4877
  signal tmp_ivl_42411 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4877
  signal tmp_ivl_42413 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4877
  signal tmp_ivl_42418 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4878
  signal tmp_ivl_42423 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4878
  signal tmp_ivl_42425 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4878
  signal tmp_ivl_42430 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4878
  signal tmp_ivl_42433 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4878
  signal tmp_ivl_42437 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4878
  signal tmp_ivl_42439 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4878
  signal tmp_ivl_42441 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4878
  signal tmp_ivl_42446 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4879
  signal tmp_ivl_4245 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3087
  signal tmp_ivl_42451 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4879
  signal tmp_ivl_42453 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4879
  signal tmp_ivl_42458 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4879
  signal tmp_ivl_42461 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4879
  signal tmp_ivl_42465 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4879
  signal tmp_ivl_42467 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4879
  signal tmp_ivl_42469 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4879
  signal tmp_ivl_4247 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3087
  signal tmp_ivl_42474 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4880
  signal tmp_ivl_42479 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4880
  signal tmp_ivl_42481 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4880
  signal tmp_ivl_42486 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4880
  signal tmp_ivl_42489 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4880
  signal tmp_ivl_42493 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4880
  signal tmp_ivl_42495 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4880
  signal tmp_ivl_42497 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4880
  signal tmp_ivl_42502 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4881
  signal tmp_ivl_42507 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4881
  signal tmp_ivl_42509 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4881
  signal tmp_ivl_42514 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4881
  signal tmp_ivl_42517 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4881
  signal tmp_ivl_42521 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4881
  signal tmp_ivl_42523 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4881
  signal tmp_ivl_42525 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4881
  signal tmp_ivl_4253 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3088
  signal tmp_ivl_42530 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4882
  signal tmp_ivl_42535 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4882
  signal tmp_ivl_42537 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4882
  signal tmp_ivl_42542 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4882
  signal tmp_ivl_42545 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4882
  signal tmp_ivl_42549 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4882
  signal tmp_ivl_4255 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3088
  signal tmp_ivl_42551 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4882
  signal tmp_ivl_42553 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4882
  signal tmp_ivl_42558 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4883
  signal tmp_ivl_4256 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3088
  signal tmp_ivl_42563 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4883
  signal tmp_ivl_42565 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4883
  signal tmp_ivl_42570 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4883
  signal tmp_ivl_42573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4883
  signal tmp_ivl_42577 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4883
  signal tmp_ivl_42579 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4883
  signal tmp_ivl_42581 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4883
  signal tmp_ivl_42586 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4884
  signal tmp_ivl_42591 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4884
  signal tmp_ivl_42593 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4884
  signal tmp_ivl_42598 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4884
  signal tmp_ivl_426 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2954
  signal tmp_ivl_42601 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4884
  signal tmp_ivl_42605 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4884
  signal tmp_ivl_42607 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4884
  signal tmp_ivl_42609 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4884
  signal tmp_ivl_4261 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3088
  signal tmp_ivl_42614 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4885
  signal tmp_ivl_42619 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4885
  signal tmp_ivl_42621 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4885
  signal tmp_ivl_42626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4885
  signal tmp_ivl_42629 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4885
  signal tmp_ivl_42633 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4885
  signal tmp_ivl_42635 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4885
  signal tmp_ivl_42637 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4885
  signal tmp_ivl_4264 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3088
  signal tmp_ivl_42642 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4886
  signal tmp_ivl_42647 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4886
  signal tmp_ivl_42649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4886
  signal tmp_ivl_42654 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4886
  signal tmp_ivl_42657 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4886
  signal tmp_ivl_4266 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3088
  signal tmp_ivl_42661 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4886
  signal tmp_ivl_42663 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4886
  signal tmp_ivl_42665 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4886
  signal tmp_ivl_4267 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3088
  signal tmp_ivl_42670 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4887
  signal tmp_ivl_42675 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4887
  signal tmp_ivl_42677 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4887
  signal tmp_ivl_42682 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4887
  signal tmp_ivl_42685 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4887
  signal tmp_ivl_42689 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4887
  signal tmp_ivl_42691 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4887
  signal tmp_ivl_42693 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4887
  signal tmp_ivl_42698 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4888
  signal tmp_ivl_42703 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4888
  signal tmp_ivl_42705 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4888
  signal tmp_ivl_42710 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4888
  signal tmp_ivl_42713 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4888
  signal tmp_ivl_42717 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4888
  signal tmp_ivl_42719 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4888
  signal tmp_ivl_4272 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3088
  signal tmp_ivl_42721 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4888
  signal tmp_ivl_42726 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4889
  signal tmp_ivl_42731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4889
  signal tmp_ivl_42733 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4889
  signal tmp_ivl_42738 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4889
  signal tmp_ivl_4274 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3088
  signal tmp_ivl_42741 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4889
  signal tmp_ivl_42745 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4889
  signal tmp_ivl_42747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4889
  signal tmp_ivl_42749 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4889
  signal tmp_ivl_42754 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4890
  signal tmp_ivl_42759 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4890
  signal tmp_ivl_42761 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4890
  signal tmp_ivl_42766 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4890
  signal tmp_ivl_42769 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4890
  signal tmp_ivl_42773 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4890
  signal tmp_ivl_42775 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4890
  signal tmp_ivl_42777 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4890
  signal tmp_ivl_42782 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4891
  signal tmp_ivl_42787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4891
  signal tmp_ivl_42789 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4891
  signal tmp_ivl_42794 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4891
  signal tmp_ivl_42797 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4891
  signal tmp_ivl_428 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2954
  signal tmp_ivl_4280 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3089
  signal tmp_ivl_42801 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4891
  signal tmp_ivl_42803 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4891
  signal tmp_ivl_42805 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4891
  signal tmp_ivl_42810 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4892
  signal tmp_ivl_42815 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4892
  signal tmp_ivl_42817 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4892
  signal tmp_ivl_4282 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3089
  signal tmp_ivl_42822 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4892
  signal tmp_ivl_42825 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4892
  signal tmp_ivl_42829 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4892
  signal tmp_ivl_4283 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3089
  signal tmp_ivl_42831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4892
  signal tmp_ivl_42833 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4892
  signal tmp_ivl_42838 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4893
  signal tmp_ivl_42843 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4893
  signal tmp_ivl_42845 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4893
  signal tmp_ivl_42850 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4893
  signal tmp_ivl_42853 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4893
  signal tmp_ivl_42857 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4893
  signal tmp_ivl_42859 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4893
  signal tmp_ivl_42861 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4893
  signal tmp_ivl_42866 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4894
  signal tmp_ivl_42871 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4894
  signal tmp_ivl_42873 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4894
  signal tmp_ivl_42878 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4894
  signal tmp_ivl_4288 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3089
  signal tmp_ivl_42881 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4894
  signal tmp_ivl_42885 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4894
  signal tmp_ivl_42887 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4894
  signal tmp_ivl_42889 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4894
  signal tmp_ivl_42894 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4895
  signal tmp_ivl_42899 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4895
  signal tmp_ivl_42901 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4895
  signal tmp_ivl_42906 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4895
  signal tmp_ivl_42909 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4895
  signal tmp_ivl_4291 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3089
  signal tmp_ivl_42913 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4895
  signal tmp_ivl_42915 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4895
  signal tmp_ivl_42917 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4895
  signal tmp_ivl_42922 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4896
  signal tmp_ivl_42927 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4896
  signal tmp_ivl_42929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4896
  signal tmp_ivl_4293 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3089
  signal tmp_ivl_42934 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4896
  signal tmp_ivl_42937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4896
  signal tmp_ivl_4294 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3089
  signal tmp_ivl_42941 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4896
  signal tmp_ivl_42943 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4896
  signal tmp_ivl_42945 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4896
  signal tmp_ivl_42950 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4897
  signal tmp_ivl_42955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4897
  signal tmp_ivl_42957 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4897
  signal tmp_ivl_42962 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4897
  signal tmp_ivl_42965 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4897
  signal tmp_ivl_42969 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4897
  signal tmp_ivl_42971 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4897
  signal tmp_ivl_42973 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4897
  signal tmp_ivl_42978 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4898
  signal tmp_ivl_42983 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4898
  signal tmp_ivl_42985 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4898
  signal tmp_ivl_4299 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3089
  signal tmp_ivl_42990 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4898
  signal tmp_ivl_42993 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4898
  signal tmp_ivl_42997 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4898
  signal tmp_ivl_42999 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4898
  signal tmp_ivl_43 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2941
  signal tmp_ivl_430 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2954
  signal tmp_ivl_43001 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4898
  signal tmp_ivl_43006 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4899
  signal tmp_ivl_4301 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3089
  signal tmp_ivl_43011 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4899
  signal tmp_ivl_43013 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4899
  signal tmp_ivl_43018 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4899
  signal tmp_ivl_43021 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4899
  signal tmp_ivl_43025 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4899
  signal tmp_ivl_43027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4899
  signal tmp_ivl_43029 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4899
  signal tmp_ivl_43034 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4900
  signal tmp_ivl_43039 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4900
  signal tmp_ivl_43041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4900
  signal tmp_ivl_43046 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4900
  signal tmp_ivl_43049 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4900
  signal tmp_ivl_43053 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4900
  signal tmp_ivl_43055 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4900
  signal tmp_ivl_43057 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4900
  signal tmp_ivl_43062 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4901
  signal tmp_ivl_43067 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4901
  signal tmp_ivl_43069 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4901
  signal tmp_ivl_4307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3090
  signal tmp_ivl_43074 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4901
  signal tmp_ivl_43077 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4901
  signal tmp_ivl_43081 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4901
  signal tmp_ivl_43083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4901
  signal tmp_ivl_43085 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4901
  signal tmp_ivl_4309 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3090
  signal tmp_ivl_43090 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4902
  signal tmp_ivl_43095 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4902
  signal tmp_ivl_43097 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4902
  signal tmp_ivl_4310 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3090
  signal tmp_ivl_43102 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4902
  signal tmp_ivl_43105 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4902
  signal tmp_ivl_43109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4902
  signal tmp_ivl_43111 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4902
  signal tmp_ivl_43113 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4902
  signal tmp_ivl_43118 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4903
  signal tmp_ivl_43123 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4903
  signal tmp_ivl_43125 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4903
  signal tmp_ivl_43130 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4903
  signal tmp_ivl_43133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4903
  signal tmp_ivl_43137 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4903
  signal tmp_ivl_43139 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4903
  signal tmp_ivl_43141 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4903
  signal tmp_ivl_43146 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4904
  signal tmp_ivl_4315 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3090
  signal tmp_ivl_43151 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4904
  signal tmp_ivl_43153 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4904
  signal tmp_ivl_43158 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4904
  signal tmp_ivl_43161 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4904
  signal tmp_ivl_43165 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4904
  signal tmp_ivl_43167 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4904
  signal tmp_ivl_43169 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4904
  signal tmp_ivl_43174 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4905
  signal tmp_ivl_43179 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4905
  signal tmp_ivl_4318 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3090
  signal tmp_ivl_43181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4905
  signal tmp_ivl_43186 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4905
  signal tmp_ivl_43189 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4905
  signal tmp_ivl_43193 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4905
  signal tmp_ivl_43195 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4905
  signal tmp_ivl_43197 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4905
  signal tmp_ivl_4320 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3090
  signal tmp_ivl_43202 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4906
  signal tmp_ivl_43207 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4906
  signal tmp_ivl_43209 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4906
  signal tmp_ivl_4321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3090
  signal tmp_ivl_43214 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4906
  signal tmp_ivl_43217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4906
  signal tmp_ivl_43221 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4906
  signal tmp_ivl_43223 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4906
  signal tmp_ivl_43225 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4906
  signal tmp_ivl_43230 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4907
  signal tmp_ivl_43235 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4907
  signal tmp_ivl_43237 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4907
  signal tmp_ivl_43242 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4907
  signal tmp_ivl_43245 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4907
  signal tmp_ivl_43249 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4907
  signal tmp_ivl_43251 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4907
  signal tmp_ivl_43253 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4907
  signal tmp_ivl_43258 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4908
  signal tmp_ivl_4326 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3090
  signal tmp_ivl_43263 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4908
  signal tmp_ivl_43265 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4908
  signal tmp_ivl_43270 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4908
  signal tmp_ivl_43273 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4908
  signal tmp_ivl_43277 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4908
  signal tmp_ivl_43279 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4908
  signal tmp_ivl_4328 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3090
  signal tmp_ivl_43281 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4908
  signal tmp_ivl_43286 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4909
  signal tmp_ivl_43291 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4909
  signal tmp_ivl_43293 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4909
  signal tmp_ivl_43298 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4909
  signal tmp_ivl_43301 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4909
  signal tmp_ivl_43305 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4909
  signal tmp_ivl_43307 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4909
  signal tmp_ivl_43309 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4909
  signal tmp_ivl_43314 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4910
  signal tmp_ivl_43319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4910
  signal tmp_ivl_43321 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4910
  signal tmp_ivl_43326 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4910
  signal tmp_ivl_43329 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4910
  signal tmp_ivl_43333 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4910
  signal tmp_ivl_43335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4910
  signal tmp_ivl_43337 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4910
  signal tmp_ivl_4334 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3091
  signal tmp_ivl_43342 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4911
  signal tmp_ivl_43347 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4911
  signal tmp_ivl_43349 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4911
  signal tmp_ivl_43354 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4911
  signal tmp_ivl_43357 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4911
  signal tmp_ivl_4336 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3091
  signal tmp_ivl_43361 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4911
  signal tmp_ivl_43363 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4911
  signal tmp_ivl_43365 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4911
  signal tmp_ivl_4337 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3091
  signal tmp_ivl_43370 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4912
  signal tmp_ivl_43375 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4912
  signal tmp_ivl_43377 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4912
  signal tmp_ivl_43382 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4912
  signal tmp_ivl_43385 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4912
  signal tmp_ivl_43389 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4912
  signal tmp_ivl_43391 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4912
  signal tmp_ivl_43393 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4912
  signal tmp_ivl_43398 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4913
  signal tmp_ivl_43403 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4913
  signal tmp_ivl_43405 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4913
  signal tmp_ivl_43410 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4913
  signal tmp_ivl_43413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4913
  signal tmp_ivl_43417 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4913
  signal tmp_ivl_43419 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4913
  signal tmp_ivl_4342 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3091
  signal tmp_ivl_43421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4913
  signal tmp_ivl_43426 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4914
  signal tmp_ivl_43431 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4914
  signal tmp_ivl_43433 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4914
  signal tmp_ivl_43438 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4914
  signal tmp_ivl_43441 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4914
  signal tmp_ivl_43445 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4914
  signal tmp_ivl_43447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4914
  signal tmp_ivl_43449 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4914
  signal tmp_ivl_4345 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3091
  signal tmp_ivl_43454 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4915
  signal tmp_ivl_43459 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4915
  signal tmp_ivl_43461 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4915
  signal tmp_ivl_43466 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4915
  signal tmp_ivl_43469 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4915
  signal tmp_ivl_4347 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3091
  signal tmp_ivl_43473 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4915
  signal tmp_ivl_43475 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4915
  signal tmp_ivl_43477 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4915
  signal tmp_ivl_4348 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3091
  signal tmp_ivl_43482 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4916
  signal tmp_ivl_43487 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4916
  signal tmp_ivl_43489 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4916
  signal tmp_ivl_43494 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4916
  signal tmp_ivl_43497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4916
  signal tmp_ivl_43501 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4916
  signal tmp_ivl_43503 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4916
  signal tmp_ivl_43505 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4916
  signal tmp_ivl_43510 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4917
  signal tmp_ivl_43515 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4917
  signal tmp_ivl_43517 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4917
  signal tmp_ivl_43522 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4917
  signal tmp_ivl_43525 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4917
  signal tmp_ivl_43529 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4917
  signal tmp_ivl_4353 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3091
  signal tmp_ivl_43531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4917
  signal tmp_ivl_43533 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4917
  signal tmp_ivl_43538 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4918
  signal tmp_ivl_43543 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4918
  signal tmp_ivl_43545 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4918
  signal tmp_ivl_4355 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3091
  signal tmp_ivl_43550 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4918
  signal tmp_ivl_43553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4918
  signal tmp_ivl_43557 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4918
  signal tmp_ivl_43559 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4918
  signal tmp_ivl_43561 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4918
  signal tmp_ivl_43566 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4919
  signal tmp_ivl_43571 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4919
  signal tmp_ivl_43573 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4919
  signal tmp_ivl_43578 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4919
  signal tmp_ivl_43581 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4919
  signal tmp_ivl_43585 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4919
  signal tmp_ivl_43587 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4919
  signal tmp_ivl_43589 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4919
  signal tmp_ivl_43594 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4920
  signal tmp_ivl_43599 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4920
  signal tmp_ivl_436 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2955
  signal tmp_ivl_43601 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4920
  signal tmp_ivl_43606 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4920
  signal tmp_ivl_43609 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4920
  signal tmp_ivl_4361 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3092
  signal tmp_ivl_43613 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4920
  signal tmp_ivl_43615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4920
  signal tmp_ivl_43617 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4920
  signal tmp_ivl_43622 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4921
  signal tmp_ivl_43627 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4921
  signal tmp_ivl_43629 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4921
  signal tmp_ivl_4363 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3092
  signal tmp_ivl_43634 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4921
  signal tmp_ivl_43637 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4921
  signal tmp_ivl_4364 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3092
  signal tmp_ivl_43641 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4921
  signal tmp_ivl_43643 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4921
  signal tmp_ivl_43645 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4921
  signal tmp_ivl_43650 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4922
  signal tmp_ivl_43655 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4922
  signal tmp_ivl_43657 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4922
  signal tmp_ivl_43662 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4922
  signal tmp_ivl_43665 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4922
  signal tmp_ivl_43669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4922
  signal tmp_ivl_43671 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4922
  signal tmp_ivl_43673 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4922
  signal tmp_ivl_43678 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4923
  signal tmp_ivl_43683 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4923
  signal tmp_ivl_43685 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4923
  signal tmp_ivl_4369 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3092
  signal tmp_ivl_43690 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4923
  signal tmp_ivl_43693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4923
  signal tmp_ivl_43697 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4923
  signal tmp_ivl_43699 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4923
  signal tmp_ivl_43701 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4923
  signal tmp_ivl_43706 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4924
  signal tmp_ivl_43711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4924
  signal tmp_ivl_43714 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4924
  signal tmp_ivl_43715 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4924
  signal tmp_ivl_4372 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3092
  signal tmp_ivl_43720 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4924
  signal tmp_ivl_43723 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4924
  signal tmp_ivl_43727 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4924
  signal tmp_ivl_43729 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4924
  signal tmp_ivl_43731 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4924
  signal tmp_ivl_43736 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4925
  signal tmp_ivl_4374 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3092
  signal tmp_ivl_43741 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4925
  signal tmp_ivl_43744 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4925
  signal tmp_ivl_43745 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4925
  signal tmp_ivl_4375 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3092
  signal tmp_ivl_43750 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4925
  signal tmp_ivl_43753 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4925
  signal tmp_ivl_43757 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4925
  signal tmp_ivl_43759 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4925
  signal tmp_ivl_43761 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4925
  signal tmp_ivl_43766 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4926
  signal tmp_ivl_43771 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4926
  signal tmp_ivl_43774 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4926
  signal tmp_ivl_43775 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4926
  signal tmp_ivl_43780 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4926
  signal tmp_ivl_43783 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4926
  signal tmp_ivl_43787 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4926
  signal tmp_ivl_43789 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4926
  signal tmp_ivl_43791 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4926
  signal tmp_ivl_43796 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4927
  signal tmp_ivl_438 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2955
  signal tmp_ivl_4380 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3092
  signal tmp_ivl_43801 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4927
  signal tmp_ivl_43804 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4927
  signal tmp_ivl_43805 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4927
  signal tmp_ivl_43810 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4927
  signal tmp_ivl_43813 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4927
  signal tmp_ivl_43817 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4927
  signal tmp_ivl_43819 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4927
  signal tmp_ivl_4382 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3092
  signal tmp_ivl_43821 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4927
  signal tmp_ivl_43826 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4928
  signal tmp_ivl_43831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4928
  signal tmp_ivl_43834 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4928
  signal tmp_ivl_43835 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4928
  signal tmp_ivl_43840 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4928
  signal tmp_ivl_43843 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4928
  signal tmp_ivl_43847 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4928
  signal tmp_ivl_43849 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4928
  signal tmp_ivl_43851 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4928
  signal tmp_ivl_43856 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4929
  signal tmp_ivl_43861 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4929
  signal tmp_ivl_43864 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4929
  signal tmp_ivl_43865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4929
  signal tmp_ivl_43870 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4929
  signal tmp_ivl_43873 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4929
  signal tmp_ivl_43877 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4929
  signal tmp_ivl_43879 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4929
  signal tmp_ivl_4388 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3093
  signal tmp_ivl_43881 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4929
  signal tmp_ivl_43886 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4930
  signal tmp_ivl_43891 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4930
  signal tmp_ivl_43894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4930
  signal tmp_ivl_43895 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4930
  signal tmp_ivl_439 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2955
  signal tmp_ivl_4390 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3093
  signal tmp_ivl_43900 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4930
  signal tmp_ivl_43903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4930
  signal tmp_ivl_43907 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4930
  signal tmp_ivl_43909 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4930
  signal tmp_ivl_4391 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3093
  signal tmp_ivl_43911 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4930
  signal tmp_ivl_43916 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4931
  signal tmp_ivl_43921 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4931
  signal tmp_ivl_43924 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4931
  signal tmp_ivl_43925 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4931
  signal tmp_ivl_43930 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4931
  signal tmp_ivl_43933 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4931
  signal tmp_ivl_43937 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4931
  signal tmp_ivl_43939 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4931
  signal tmp_ivl_43941 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4931
  signal tmp_ivl_43946 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4932
  signal tmp_ivl_43951 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4932
  signal tmp_ivl_43954 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4932
  signal tmp_ivl_43955 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4932
  signal tmp_ivl_4396 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3093
  signal tmp_ivl_43960 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4932
  signal tmp_ivl_43963 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4932
  signal tmp_ivl_43967 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4932
  signal tmp_ivl_43969 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4932
  signal tmp_ivl_43971 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4932
  signal tmp_ivl_43976 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4933
  signal tmp_ivl_43981 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4933
  signal tmp_ivl_43984 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4933
  signal tmp_ivl_43985 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4933
  signal tmp_ivl_4399 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3093
  signal tmp_ivl_43990 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4933
  signal tmp_ivl_43993 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4933
  signal tmp_ivl_43997 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4933
  signal tmp_ivl_43999 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4933
  signal tmp_ivl_44 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2941
  signal tmp_ivl_44001 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4933
  signal tmp_ivl_44006 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4934
  signal tmp_ivl_4401 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3093
  signal tmp_ivl_44011 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4934
  signal tmp_ivl_44014 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4934
  signal tmp_ivl_44015 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4934
  signal tmp_ivl_4402 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3093
  signal tmp_ivl_44020 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4934
  signal tmp_ivl_44023 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4934
  signal tmp_ivl_44027 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4934
  signal tmp_ivl_44029 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4934
  signal tmp_ivl_44031 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4934
  signal tmp_ivl_44036 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4935
  signal tmp_ivl_44041 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4935
  signal tmp_ivl_44044 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4935
  signal tmp_ivl_44045 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4935
  signal tmp_ivl_44050 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4935
  signal tmp_ivl_44053 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4935
  signal tmp_ivl_44057 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4935
  signal tmp_ivl_44059 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4935
  signal tmp_ivl_44061 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4935
  signal tmp_ivl_44066 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4936
  signal tmp_ivl_4407 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3093
  signal tmp_ivl_44071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4936
  signal tmp_ivl_44074 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4936
  signal tmp_ivl_44075 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4936
  signal tmp_ivl_44080 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4936
  signal tmp_ivl_44083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4936
  signal tmp_ivl_44087 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4936
  signal tmp_ivl_44089 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4936
  signal tmp_ivl_4409 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3093
  signal tmp_ivl_44091 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4936
  signal tmp_ivl_44096 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4937
  signal tmp_ivl_44101 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4937
  signal tmp_ivl_44104 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4937
  signal tmp_ivl_44105 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4937
  signal tmp_ivl_44110 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4937
  signal tmp_ivl_44113 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4937
  signal tmp_ivl_44117 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4937
  signal tmp_ivl_44119 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4937
  signal tmp_ivl_44121 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4937
  signal tmp_ivl_44126 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4938
  signal tmp_ivl_44131 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4938
  signal tmp_ivl_44134 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4938
  signal tmp_ivl_44135 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4938
  signal tmp_ivl_44140 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4938
  signal tmp_ivl_44143 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4938
  signal tmp_ivl_44147 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4938
  signal tmp_ivl_44149 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4938
  signal tmp_ivl_4415 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3094
  signal tmp_ivl_44151 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4938
  signal tmp_ivl_44156 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4939
  signal tmp_ivl_44161 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4939
  signal tmp_ivl_44164 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4939
  signal tmp_ivl_44165 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4939
  signal tmp_ivl_4417 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3094
  signal tmp_ivl_44170 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4939
  signal tmp_ivl_44173 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4939
  signal tmp_ivl_44177 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4939
  signal tmp_ivl_44179 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4939
  signal tmp_ivl_4418 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3094
  signal tmp_ivl_44181 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4939
  signal tmp_ivl_44186 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4940
  signal tmp_ivl_44191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4940
  signal tmp_ivl_44194 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4940
  signal tmp_ivl_44195 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4940
  signal tmp_ivl_44200 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4940
  signal tmp_ivl_44203 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4940
  signal tmp_ivl_44207 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4940
  signal tmp_ivl_44209 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4940
  signal tmp_ivl_44211 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4940
  signal tmp_ivl_44216 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4941
  signal tmp_ivl_44221 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4941
  signal tmp_ivl_44224 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4941
  signal tmp_ivl_44225 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4941
  signal tmp_ivl_4423 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3094
  signal tmp_ivl_44230 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4941
  signal tmp_ivl_44233 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4941
  signal tmp_ivl_44237 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4941
  signal tmp_ivl_44239 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4941
  signal tmp_ivl_44241 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4941
  signal tmp_ivl_44246 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4942
  signal tmp_ivl_44251 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4942
  signal tmp_ivl_44254 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4942
  signal tmp_ivl_44255 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4942
  signal tmp_ivl_4426 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3094
  signal tmp_ivl_44260 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4942
  signal tmp_ivl_44263 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4942
  signal tmp_ivl_44267 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4942
  signal tmp_ivl_44269 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4942
  signal tmp_ivl_44271 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4942
  signal tmp_ivl_44276 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4943
  signal tmp_ivl_4428 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3094
  signal tmp_ivl_44281 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4943
  signal tmp_ivl_44284 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4943
  signal tmp_ivl_44285 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4943
  signal tmp_ivl_4429 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3094
  signal tmp_ivl_44290 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4943
  signal tmp_ivl_44293 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4943
  signal tmp_ivl_44297 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4943
  signal tmp_ivl_44299 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4943
  signal tmp_ivl_44301 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4943
  signal tmp_ivl_44306 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4944
  signal tmp_ivl_44311 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4944
  signal tmp_ivl_44314 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4944
  signal tmp_ivl_44315 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4944
  signal tmp_ivl_44320 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4944
  signal tmp_ivl_44323 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4944
  signal tmp_ivl_44327 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4944
  signal tmp_ivl_44329 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4944
  signal tmp_ivl_44331 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4944
  signal tmp_ivl_44336 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4945
  signal tmp_ivl_4434 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3094
  signal tmp_ivl_44341 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4945
  signal tmp_ivl_44344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4945
  signal tmp_ivl_44345 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4945
  signal tmp_ivl_44350 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4945
  signal tmp_ivl_44353 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4945
  signal tmp_ivl_44357 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4945
  signal tmp_ivl_44359 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4945
  signal tmp_ivl_4436 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3094
  signal tmp_ivl_44361 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4945
  signal tmp_ivl_44366 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4946
  signal tmp_ivl_44371 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4946
  signal tmp_ivl_44374 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4946
  signal tmp_ivl_44375 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4946
  signal tmp_ivl_44380 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4946
  signal tmp_ivl_44383 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4946
  signal tmp_ivl_44387 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4946
  signal tmp_ivl_44389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4946
  signal tmp_ivl_44391 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4946
  signal tmp_ivl_44396 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4947
  signal tmp_ivl_444 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2955
  signal tmp_ivl_44401 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4947
  signal tmp_ivl_44404 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4947
  signal tmp_ivl_44405 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4947
  signal tmp_ivl_44410 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4947
  signal tmp_ivl_44413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4947
  signal tmp_ivl_44417 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4947
  signal tmp_ivl_44419 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4947
  signal tmp_ivl_4442 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3095
  signal tmp_ivl_44421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4947
  signal tmp_ivl_44426 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4948
  signal tmp_ivl_44431 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4948
  signal tmp_ivl_44434 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4948
  signal tmp_ivl_44435 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4948
  signal tmp_ivl_4444 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3095
  signal tmp_ivl_44440 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4948
  signal tmp_ivl_44443 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4948
  signal tmp_ivl_44447 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4948
  signal tmp_ivl_44449 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4948
  signal tmp_ivl_4445 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3095
  signal tmp_ivl_44451 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4948
  signal tmp_ivl_44456 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4949
  signal tmp_ivl_44461 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4949
  signal tmp_ivl_44464 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4949
  signal tmp_ivl_44465 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4949
  signal tmp_ivl_44470 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4949
  signal tmp_ivl_44473 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4949
  signal tmp_ivl_44477 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4949
  signal tmp_ivl_44479 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4949
  signal tmp_ivl_44481 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4949
  signal tmp_ivl_4450 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3095
  signal tmp_ivl_4453 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3095
  signal tmp_ivl_4455 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3095
  signal tmp_ivl_4456 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3095
  signal tmp_ivl_4461 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3095
  signal tmp_ivl_4463 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3095
  signal tmp_ivl_4469 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3096
  signal tmp_ivl_447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2955
  signal tmp_ivl_4471 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3096
  signal tmp_ivl_4472 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3096
  signal tmp_ivl_4477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3096
  signal tmp_ivl_4480 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3096
  signal tmp_ivl_4482 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3096
  signal tmp_ivl_4483 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3096
  signal tmp_ivl_4488 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3096
  signal tmp_ivl_449 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2955
  signal tmp_ivl_4490 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3096
  signal tmp_ivl_4496 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3097
  signal tmp_ivl_4498 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3097
  signal tmp_ivl_4499 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3097
  signal tmp_ivl_450 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2955
  signal tmp_ivl_4504 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3097
  signal tmp_ivl_4507 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3097
  signal tmp_ivl_4509 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3097
  signal tmp_ivl_4510 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3097
  signal tmp_ivl_4515 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3097
  signal tmp_ivl_4517 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3097
  signal tmp_ivl_4523 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3098
  signal tmp_ivl_4525 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3098
  signal tmp_ivl_4526 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3098
  signal tmp_ivl_4531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3098
  signal tmp_ivl_4534 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3098
  signal tmp_ivl_4536 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3098
  signal tmp_ivl_4537 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3098
  signal tmp_ivl_4542 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3098
  signal tmp_ivl_4544 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3098
  signal tmp_ivl_455 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2955
  signal tmp_ivl_4550 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3099
  signal tmp_ivl_4552 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3099
  signal tmp_ivl_4553 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3099
  signal tmp_ivl_4558 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3099
  signal tmp_ivl_4561 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3099
  signal tmp_ivl_4563 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3099
  signal tmp_ivl_4564 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3099
  signal tmp_ivl_4569 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3099
  signal tmp_ivl_457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2955
  signal tmp_ivl_4571 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3099
  signal tmp_ivl_4577 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3100
  signal tmp_ivl_4579 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3100
  signal tmp_ivl_4580 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3100
  signal tmp_ivl_4585 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3100
  signal tmp_ivl_4588 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3100
  signal tmp_ivl_459 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2955
  signal tmp_ivl_4590 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3100
  signal tmp_ivl_4591 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3100
  signal tmp_ivl_4596 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3100
  signal tmp_ivl_4598 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3100
  signal tmp_ivl_4604 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3101
  signal tmp_ivl_4606 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3101
  signal tmp_ivl_4607 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3101
  signal tmp_ivl_4612 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3101
  signal tmp_ivl_4615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3101
  signal tmp_ivl_4617 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3101
  signal tmp_ivl_4618 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3101
  signal tmp_ivl_4623 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3101
  signal tmp_ivl_4625 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3101
  signal tmp_ivl_4631 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3102
  signal tmp_ivl_4633 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3102
  signal tmp_ivl_4634 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3102
  signal tmp_ivl_4639 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3102
  signal tmp_ivl_4642 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3102
  signal tmp_ivl_4644 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3102
  signal tmp_ivl_4645 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3102
  signal tmp_ivl_465 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2956
  signal tmp_ivl_4650 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3102
  signal tmp_ivl_4652 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3102
  signal tmp_ivl_4658 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3103
  signal tmp_ivl_4660 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3103
  signal tmp_ivl_4661 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3103
  signal tmp_ivl_4666 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3103
  signal tmp_ivl_4669 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3103
  signal tmp_ivl_467 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2956
  signal tmp_ivl_4671 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3103
  signal tmp_ivl_4672 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3103
  signal tmp_ivl_4677 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3103
  signal tmp_ivl_4679 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3103
  signal tmp_ivl_468 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2956
  signal tmp_ivl_4685 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3104
  signal tmp_ivl_4687 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3104
  signal tmp_ivl_4688 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3104
  signal tmp_ivl_4693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3104
  signal tmp_ivl_4696 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3104
  signal tmp_ivl_4698 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3104
  signal tmp_ivl_4699 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3104
  signal tmp_ivl_4704 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3104
  signal tmp_ivl_4706 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3104
  signal tmp_ivl_4712 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3105
  signal tmp_ivl_4714 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3105
  signal tmp_ivl_4715 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3105
  signal tmp_ivl_4720 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3105
  signal tmp_ivl_4723 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3105
  signal tmp_ivl_4725 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3105
  signal tmp_ivl_4726 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3105
  signal tmp_ivl_473 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2956
  signal tmp_ivl_4731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3105
  signal tmp_ivl_4733 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3105
  signal tmp_ivl_4739 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3106
  signal tmp_ivl_4741 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3106
  signal tmp_ivl_4742 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3106
  signal tmp_ivl_4747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3106
  signal tmp_ivl_4750 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3106
  signal tmp_ivl_4752 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3106
  signal tmp_ivl_4753 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3106
  signal tmp_ivl_4758 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3106
  signal tmp_ivl_476 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2956
  signal tmp_ivl_4760 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3106
  signal tmp_ivl_4766 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3107
  signal tmp_ivl_4768 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3107
  signal tmp_ivl_4769 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3107
  signal tmp_ivl_4774 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3107
  signal tmp_ivl_4777 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3107
  signal tmp_ivl_4779 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3107
  signal tmp_ivl_478 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2956
  signal tmp_ivl_4780 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3107
  signal tmp_ivl_4785 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3107
  signal tmp_ivl_4787 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3107
  signal tmp_ivl_479 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2956
  signal tmp_ivl_4793 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3108
  signal tmp_ivl_4795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3108
  signal tmp_ivl_4796 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3108
  signal tmp_ivl_4801 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3108
  signal tmp_ivl_4804 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3108
  signal tmp_ivl_4806 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3108
  signal tmp_ivl_4807 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3108
  signal tmp_ivl_4812 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3108
  signal tmp_ivl_4814 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3108
  signal tmp_ivl_4820 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3109
  signal tmp_ivl_4822 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3109
  signal tmp_ivl_4823 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3109
  signal tmp_ivl_4828 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3109
  signal tmp_ivl_4831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3109
  signal tmp_ivl_4833 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3109
  signal tmp_ivl_4834 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3109
  signal tmp_ivl_4839 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3109
  signal tmp_ivl_484 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2956
  signal tmp_ivl_4841 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3109
  signal tmp_ivl_4847 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3110
  signal tmp_ivl_4849 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3110
  signal tmp_ivl_4850 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3110
  signal tmp_ivl_4855 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3110
  signal tmp_ivl_4858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3110
  signal tmp_ivl_486 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2956
  signal tmp_ivl_4860 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3110
  signal tmp_ivl_4861 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3110
  signal tmp_ivl_4866 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3110
  signal tmp_ivl_4868 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3110
  signal tmp_ivl_4874 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3111
  signal tmp_ivl_4876 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3111
  signal tmp_ivl_4877 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3111
  signal tmp_ivl_488 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2956
  signal tmp_ivl_4882 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3111
  signal tmp_ivl_4885 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3111
  signal tmp_ivl_4887 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3111
  signal tmp_ivl_4888 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3111
  signal tmp_ivl_4893 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3111
  signal tmp_ivl_4895 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3111
  signal tmp_ivl_49 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2941
  signal tmp_ivl_4901 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3112
  signal tmp_ivl_4903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3112
  signal tmp_ivl_4904 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3112
  signal tmp_ivl_4909 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3112
  signal tmp_ivl_4912 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3112
  signal tmp_ivl_4914 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3112
  signal tmp_ivl_4915 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3112
  signal tmp_ivl_4920 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3112
  signal tmp_ivl_4922 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3112
  signal tmp_ivl_4928 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3113
  signal tmp_ivl_4930 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3113
  signal tmp_ivl_4931 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3113
  signal tmp_ivl_4936 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3113
  signal tmp_ivl_4939 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3113
  signal tmp_ivl_494 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2957
  signal tmp_ivl_4941 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3113
  signal tmp_ivl_4942 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3113
  signal tmp_ivl_4947 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3113
  signal tmp_ivl_4949 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3113
  signal tmp_ivl_4955 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3114
  signal tmp_ivl_4957 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3114
  signal tmp_ivl_4958 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3114
  signal tmp_ivl_496 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2957
  signal tmp_ivl_4963 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3114
  signal tmp_ivl_4966 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3114
  signal tmp_ivl_4968 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3114
  signal tmp_ivl_4969 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3114
  signal tmp_ivl_497 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2957
  signal tmp_ivl_4974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3114
  signal tmp_ivl_4976 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3114
  signal tmp_ivl_4982 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3115
  signal tmp_ivl_4984 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3115
  signal tmp_ivl_4985 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3115
  signal tmp_ivl_4990 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3115
  signal tmp_ivl_4993 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3115
  signal tmp_ivl_4995 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3115
  signal tmp_ivl_4996 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3115
  signal tmp_ivl_5001 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3115
  signal tmp_ivl_5003 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3115
  signal tmp_ivl_5009 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3116
  signal tmp_ivl_5011 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3116
  signal tmp_ivl_5012 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3116
  signal tmp_ivl_5017 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3116
  signal tmp_ivl_502 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2957
  signal tmp_ivl_5020 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3116
  signal tmp_ivl_5022 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3116
  signal tmp_ivl_5023 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3116
  signal tmp_ivl_5028 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3116
  signal tmp_ivl_5030 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3116
  signal tmp_ivl_5036 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3117
  signal tmp_ivl_5038 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3117
  signal tmp_ivl_5039 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3117
  signal tmp_ivl_5044 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3117
  signal tmp_ivl_5047 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3117
  signal tmp_ivl_5049 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3117
  signal tmp_ivl_505 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2957
  signal tmp_ivl_5050 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3117
  signal tmp_ivl_5055 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3117
  signal tmp_ivl_5057 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3117
  signal tmp_ivl_5063 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3118
  signal tmp_ivl_5065 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3118
  signal tmp_ivl_5066 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3118
  signal tmp_ivl_507 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2957
  signal tmp_ivl_5071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3118
  signal tmp_ivl_5074 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3118
  signal tmp_ivl_5076 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3118
  signal tmp_ivl_5077 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3118
  signal tmp_ivl_508 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2957
  signal tmp_ivl_5082 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3118
  signal tmp_ivl_5084 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3118
  signal tmp_ivl_5090 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3119
  signal tmp_ivl_5092 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3119
  signal tmp_ivl_5093 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3119
  signal tmp_ivl_5098 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3119
  signal tmp_ivl_51 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2941
  signal tmp_ivl_5101 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3119
  signal tmp_ivl_5103 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3119
  signal tmp_ivl_5104 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3119
  signal tmp_ivl_5109 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3119
  signal tmp_ivl_5111 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3119
  signal tmp_ivl_5117 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3120
  signal tmp_ivl_5119 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3120
  signal tmp_ivl_5120 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3120
  signal tmp_ivl_5125 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3120
  signal tmp_ivl_5128 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3120
  signal tmp_ivl_513 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2957
  signal tmp_ivl_5130 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3120
  signal tmp_ivl_5131 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3120
  signal tmp_ivl_5136 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3120
  signal tmp_ivl_5138 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3120
  signal tmp_ivl_5144 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3121
  signal tmp_ivl_5146 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3121
  signal tmp_ivl_5147 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3121
  signal tmp_ivl_515 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2957
  signal tmp_ivl_5152 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3121
  signal tmp_ivl_5155 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3121
  signal tmp_ivl_5157 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3121
  signal tmp_ivl_5158 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3121
  signal tmp_ivl_5163 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3121
  signal tmp_ivl_5165 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3121
  signal tmp_ivl_517 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2957
  signal tmp_ivl_5171 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3122
  signal tmp_ivl_5173 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3122
  signal tmp_ivl_5174 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3122
  signal tmp_ivl_5179 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3122
  signal tmp_ivl_5182 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3122
  signal tmp_ivl_5184 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3122
  signal tmp_ivl_5185 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3122
  signal tmp_ivl_5190 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3122
  signal tmp_ivl_5192 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3122
  signal tmp_ivl_5198 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3123
  signal tmp_ivl_5200 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3123
  signal tmp_ivl_5201 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3123
  signal tmp_ivl_5206 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3123
  signal tmp_ivl_5209 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3123
  signal tmp_ivl_5211 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3123
  signal tmp_ivl_5212 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3123
  signal tmp_ivl_5217 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3123
  signal tmp_ivl_5219 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3123
  signal tmp_ivl_5225 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3124
  signal tmp_ivl_5227 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3124
  signal tmp_ivl_5228 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3124
  signal tmp_ivl_523 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2958
  signal tmp_ivl_5233 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3124
  signal tmp_ivl_5236 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3124
  signal tmp_ivl_5238 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3124
  signal tmp_ivl_5239 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3124
  signal tmp_ivl_5244 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3124
  signal tmp_ivl_5246 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3124
  signal tmp_ivl_525 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2958
  signal tmp_ivl_5252 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3125
  signal tmp_ivl_5254 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3125
  signal tmp_ivl_5255 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3125
  signal tmp_ivl_526 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2958
  signal tmp_ivl_5260 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3125
  signal tmp_ivl_5263 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3125
  signal tmp_ivl_5265 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3125
  signal tmp_ivl_5266 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3125
  signal tmp_ivl_5271 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3125
  signal tmp_ivl_5273 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3125
  signal tmp_ivl_5279 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3126
  signal tmp_ivl_5281 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3126
  signal tmp_ivl_5282 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3126
  signal tmp_ivl_5287 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3126
  signal tmp_ivl_5290 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3126
  signal tmp_ivl_5292 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3126
  signal tmp_ivl_5293 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3126
  signal tmp_ivl_5298 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3126
  signal tmp_ivl_53 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2941
  signal tmp_ivl_5300 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3126
  signal tmp_ivl_5306 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3127
  signal tmp_ivl_5308 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3127
  signal tmp_ivl_5309 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3127
  signal tmp_ivl_531 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2958
  signal tmp_ivl_5314 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3127
  signal tmp_ivl_5317 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3127
  signal tmp_ivl_5319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3127
  signal tmp_ivl_5320 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3127
  signal tmp_ivl_5325 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3127
  signal tmp_ivl_5327 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3127
  signal tmp_ivl_5333 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3128
  signal tmp_ivl_5335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3128
  signal tmp_ivl_5336 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3128
  signal tmp_ivl_534 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2958
  signal tmp_ivl_5341 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3128
  signal tmp_ivl_5344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3128
  signal tmp_ivl_5346 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3128
  signal tmp_ivl_5347 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3128
  signal tmp_ivl_5352 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3128
  signal tmp_ivl_5354 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3128
  signal tmp_ivl_536 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2958
  signal tmp_ivl_5360 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3129
  signal tmp_ivl_5362 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3129
  signal tmp_ivl_5363 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3129
  signal tmp_ivl_5368 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3129
  signal tmp_ivl_537 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2958
  signal tmp_ivl_5371 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3129
  signal tmp_ivl_5373 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3129
  signal tmp_ivl_5374 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3129
  signal tmp_ivl_5379 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3129
  signal tmp_ivl_5381 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3129
  signal tmp_ivl_5387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3130
  signal tmp_ivl_5389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3130
  signal tmp_ivl_5390 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3130
  signal tmp_ivl_5395 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3130
  signal tmp_ivl_5398 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3130
  signal tmp_ivl_5400 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3130
  signal tmp_ivl_5401 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3130
  signal tmp_ivl_5406 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3130
  signal tmp_ivl_5408 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3130
  signal tmp_ivl_5414 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3131
  signal tmp_ivl_5416 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3131
  signal tmp_ivl_5417 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3131
  signal tmp_ivl_542 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2958
  signal tmp_ivl_5422 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3131
  signal tmp_ivl_5425 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3131
  signal tmp_ivl_5427 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3131
  signal tmp_ivl_5428 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3131
  signal tmp_ivl_5433 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3131
  signal tmp_ivl_5435 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3131
  signal tmp_ivl_544 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2958
  signal tmp_ivl_5441 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3132
  signal tmp_ivl_5443 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3132
  signal tmp_ivl_5444 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3132
  signal tmp_ivl_5449 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3132
  signal tmp_ivl_5452 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3132
  signal tmp_ivl_5454 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3132
  signal tmp_ivl_5455 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3132
  signal tmp_ivl_546 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2958
  signal tmp_ivl_5460 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3132
  signal tmp_ivl_5462 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3132
  signal tmp_ivl_5468 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3133
  signal tmp_ivl_5470 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3133
  signal tmp_ivl_5471 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3133
  signal tmp_ivl_5476 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3133
  signal tmp_ivl_5479 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3133
  signal tmp_ivl_5481 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3133
  signal tmp_ivl_5482 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3133
  signal tmp_ivl_5487 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3133
  signal tmp_ivl_5489 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3133
  signal tmp_ivl_5495 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3134
  signal tmp_ivl_5497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3134
  signal tmp_ivl_5498 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3134
  signal tmp_ivl_5503 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3134
  signal tmp_ivl_5506 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3134
  signal tmp_ivl_5508 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3134
  signal tmp_ivl_5509 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3134
  signal tmp_ivl_5514 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3134
  signal tmp_ivl_5516 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3134
  signal tmp_ivl_552 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2959
  signal tmp_ivl_5522 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3135
  signal tmp_ivl_5524 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3135
  signal tmp_ivl_5525 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3135
  signal tmp_ivl_5530 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3135
  signal tmp_ivl_5533 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3135
  signal tmp_ivl_5535 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3135
  signal tmp_ivl_5536 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3135
  signal tmp_ivl_554 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2959
  signal tmp_ivl_5541 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3135
  signal tmp_ivl_5543 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3135
  signal tmp_ivl_5549 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3136
  signal tmp_ivl_555 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2959
  signal tmp_ivl_5551 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3136
  signal tmp_ivl_5552 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3136
  signal tmp_ivl_5557 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3136
  signal tmp_ivl_5560 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3136
  signal tmp_ivl_5562 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3136
  signal tmp_ivl_5563 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3136
  signal tmp_ivl_5568 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3136
  signal tmp_ivl_5570 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3136
  signal tmp_ivl_5576 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3137
  signal tmp_ivl_5578 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3137
  signal tmp_ivl_5579 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3137
  signal tmp_ivl_5584 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3137
  signal tmp_ivl_5587 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3137
  signal tmp_ivl_5589 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3137
  signal tmp_ivl_5590 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3137
  signal tmp_ivl_5595 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3137
  signal tmp_ivl_5597 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3137
  signal tmp_ivl_560 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2959
  signal tmp_ivl_5604 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3139
  signal tmp_ivl_5609 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3139
  signal tmp_ivl_5611 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3139
  signal tmp_ivl_5613 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3139
  signal tmp_ivl_5618 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3139
  signal tmp_ivl_5620 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3139
  signal tmp_ivl_5622 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3139
  signal tmp_ivl_5628 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3140
  signal tmp_ivl_563 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2959
  signal tmp_ivl_5630 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3140
  signal tmp_ivl_5631 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3140
  signal tmp_ivl_5636 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3140
  signal tmp_ivl_5639 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3140
  signal tmp_ivl_5641 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3140
  signal tmp_ivl_5642 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3140
  signal tmp_ivl_5647 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3140
  signal tmp_ivl_5649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3140
  signal tmp_ivl_565 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2959
  signal tmp_ivl_5655 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3141
  signal tmp_ivl_5657 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3141
  signal tmp_ivl_5658 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3141
  signal tmp_ivl_566 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2959
  signal tmp_ivl_5663 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3141
  signal tmp_ivl_5666 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3141
  signal tmp_ivl_5668 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3141
  signal tmp_ivl_5669 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3141
  signal tmp_ivl_5674 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3141
  signal tmp_ivl_5676 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3141
  signal tmp_ivl_5682 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3142
  signal tmp_ivl_5684 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3142
  signal tmp_ivl_5685 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3142
  signal tmp_ivl_5690 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3142
  signal tmp_ivl_5693 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3142
  signal tmp_ivl_5695 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3142
  signal tmp_ivl_5696 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3142
  signal tmp_ivl_5701 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3142
  signal tmp_ivl_5703 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3142
  signal tmp_ivl_5709 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3143
  signal tmp_ivl_571 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2959
  signal tmp_ivl_5711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3143
  signal tmp_ivl_5712 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3143
  signal tmp_ivl_5717 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3143
  signal tmp_ivl_5720 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3143
  signal tmp_ivl_5722 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3143
  signal tmp_ivl_5723 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3143
  signal tmp_ivl_5728 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3143
  signal tmp_ivl_573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2959
  signal tmp_ivl_5730 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3143
  signal tmp_ivl_5735 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3144
  signal tmp_ivl_5738 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3144
  signal tmp_ivl_5739 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3144
  signal tmp_ivl_5744 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3144
  signal tmp_ivl_5746 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3144
  signal tmp_ivl_575 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2959
  signal tmp_ivl_5751 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3144
  signal tmp_ivl_5753 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3144
  signal tmp_ivl_5759 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3145
  signal tmp_ivl_5761 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3145
  signal tmp_ivl_5762 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3145
  signal tmp_ivl_5767 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3145
  signal tmp_ivl_5770 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3145
  signal tmp_ivl_5772 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3145
  signal tmp_ivl_5773 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3145
  signal tmp_ivl_5778 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3145
  signal tmp_ivl_5780 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3145
  signal tmp_ivl_5790 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3148
  signal tmp_ivl_5792 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3148
  signal tmp_ivl_5793 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3148
  signal tmp_ivl_5798 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3148
  signal tmp_ivl_5801 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3148
  signal tmp_ivl_5803 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3148
  signal tmp_ivl_5804 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3148
  signal tmp_ivl_5809 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3148
  signal tmp_ivl_581 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2960
  signal tmp_ivl_5811 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3148
  signal tmp_ivl_5816 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3149
  signal tmp_ivl_5818 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3149
  signal tmp_ivl_5823 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3149
  signal tmp_ivl_5825 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3149
  signal tmp_ivl_583 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2960
  signal tmp_ivl_5830 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3149
  signal tmp_ivl_5832 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3149
  signal tmp_ivl_5834 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3149
  signal tmp_ivl_584 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2960
  signal tmp_ivl_5840 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3150
  signal tmp_ivl_5842 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3150
  signal tmp_ivl_5843 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3150
  signal tmp_ivl_5848 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3150
  signal tmp_ivl_5851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3150
  signal tmp_ivl_5853 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3150
  signal tmp_ivl_5854 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3150
  signal tmp_ivl_5859 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3150
  signal tmp_ivl_5861 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3150
  signal tmp_ivl_5868 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3153
  signal tmp_ivl_5873 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3153
  signal tmp_ivl_5875 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3153
  signal tmp_ivl_5877 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3153
  signal tmp_ivl_5882 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3153
  signal tmp_ivl_5884 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3153
  signal tmp_ivl_589 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2960
  signal tmp_ivl_5893 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3156
  signal tmp_ivl_5895 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3156
  signal tmp_ivl_59 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2942
  signal tmp_ivl_5900 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3156
  signal tmp_ivl_5903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3156
  signal tmp_ivl_5905 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3156
  signal tmp_ivl_5906 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3156
  signal tmp_ivl_5911 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3156
  signal tmp_ivl_5913 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3156
  signal tmp_ivl_5919 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3157
  signal tmp_ivl_592 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2960
  signal tmp_ivl_5921 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3157
  signal tmp_ivl_5922 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3157
  signal tmp_ivl_5927 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3157
  signal tmp_ivl_5929 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3157
  signal tmp_ivl_5934 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3157
  signal tmp_ivl_5936 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3157
  signal tmp_ivl_594 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2960
  signal tmp_ivl_5941 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3158
  signal tmp_ivl_5943 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3158
  signal tmp_ivl_5948 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3158
  signal tmp_ivl_595 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2960
  signal tmp_ivl_5951 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3158
  signal tmp_ivl_5953 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3158
  signal tmp_ivl_5954 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3158
  signal tmp_ivl_5959 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3158
  signal tmp_ivl_5961 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3158
  signal tmp_ivl_5966 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3159
  signal tmp_ivl_5971 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3159
  signal tmp_ivl_5974 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3159
  signal tmp_ivl_5976 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3159
  signal tmp_ivl_5977 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3159
  signal tmp_ivl_5982 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3159
  signal tmp_ivl_5984 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3159
  signal tmp_ivl_5990 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3160
  signal tmp_ivl_5992 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3160
  signal tmp_ivl_5993 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3160
  signal tmp_ivl_5998 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3160
  signal tmp_ivl_600 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2960
  signal tmp_ivl_6001 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3160
  signal tmp_ivl_6003 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3160
  signal tmp_ivl_6004 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3160
  signal tmp_ivl_6009 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3160
  signal tmp_ivl_6011 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3160
  signal tmp_ivl_6016 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3161
  signal tmp_ivl_6018 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3161
  signal tmp_ivl_602 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2960
  signal tmp_ivl_6023 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3161
  signal tmp_ivl_6025 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3161
  signal tmp_ivl_6030 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3161
  signal tmp_ivl_6032 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3161
  signal tmp_ivl_6038 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3162
  signal tmp_ivl_604 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2960
  signal tmp_ivl_6040 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3162
  signal tmp_ivl_6041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3162
  signal tmp_ivl_6046 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3162
  signal tmp_ivl_6049 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3162
  signal tmp_ivl_6051 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3162
  signal tmp_ivl_6052 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3162
  signal tmp_ivl_6057 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3162
  signal tmp_ivl_6059 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3162
  signal tmp_ivl_6064 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3163
  signal tmp_ivl_6066 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3163
  signal tmp_ivl_6071 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3163
  signal tmp_ivl_6073 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3163
  signal tmp_ivl_6078 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3163
  signal tmp_ivl_6080 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3163
  signal tmp_ivl_6086 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3164
  signal tmp_ivl_6093 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3165
  signal tmp_ivl_61 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2942
  signal tmp_ivl_610 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2961
  signal tmp_ivl_6100 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3166
  signal tmp_ivl_6107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3167
  signal tmp_ivl_6114 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3168
  signal tmp_ivl_612 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2961
  signal tmp_ivl_6121 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3169
  signal tmp_ivl_6128 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3170
  signal tmp_ivl_613 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2961
  signal tmp_ivl_6135 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3171
  signal tmp_ivl_6142 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3172
  signal tmp_ivl_6149 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3173
  signal tmp_ivl_6156 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3174
  signal tmp_ivl_6163 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3175
  signal tmp_ivl_6170 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3176
  signal tmp_ivl_6177 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3177
  signal tmp_ivl_618 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2961
  signal tmp_ivl_6184 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3178
  signal tmp_ivl_6191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3179
  signal tmp_ivl_6198 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3180
  signal tmp_ivl_62 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2942
  signal tmp_ivl_6205 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3181
  signal tmp_ivl_621 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2961
  signal tmp_ivl_6212 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3182
  signal tmp_ivl_6219 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3183
  signal tmp_ivl_6226 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3184
  signal tmp_ivl_623 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2961
  signal tmp_ivl_6233 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3185
  signal tmp_ivl_624 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2961
  signal tmp_ivl_6240 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3186
  signal tmp_ivl_6247 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3187
  signal tmp_ivl_6254 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3188
  signal tmp_ivl_6261 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3189
  signal tmp_ivl_6268 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3190
  signal tmp_ivl_6275 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3191
  signal tmp_ivl_6282 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3192
  signal tmp_ivl_6289 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3193
  signal tmp_ivl_629 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2961
  signal tmp_ivl_6296 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3194
  signal tmp_ivl_6303 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3195
  signal tmp_ivl_631 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2961
  signal tmp_ivl_6310 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3196
  signal tmp_ivl_6317 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3197
  signal tmp_ivl_6324 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3198
  signal tmp_ivl_633 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2961
  signal tmp_ivl_6331 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3199
  signal tmp_ivl_6338 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3200
  signal tmp_ivl_6345 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3201
  signal tmp_ivl_6352 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3202
  signal tmp_ivl_6359 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3203
  signal tmp_ivl_6366 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3204
  signal tmp_ivl_6373 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3205
  signal tmp_ivl_6380 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3206
  signal tmp_ivl_6387 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3207
  signal tmp_ivl_639 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2962
  signal tmp_ivl_6394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3208
  signal tmp_ivl_6401 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3209
  signal tmp_ivl_6408 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3210
  signal tmp_ivl_641 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2962
  signal tmp_ivl_6415 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3211
  signal tmp_ivl_642 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2962
  signal tmp_ivl_6422 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3212
  signal tmp_ivl_6429 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3213
  signal tmp_ivl_6436 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3214
  signal tmp_ivl_6443 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3215
  signal tmp_ivl_6450 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3216
  signal tmp_ivl_6457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3217
  signal tmp_ivl_6464 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3218
  signal tmp_ivl_647 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2962
  signal tmp_ivl_6471 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3219
  signal tmp_ivl_6478 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3220
  signal tmp_ivl_6485 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3221
  signal tmp_ivl_6492 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3222
  signal tmp_ivl_6499 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3223
  signal tmp_ivl_650 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2962
  signal tmp_ivl_6506 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3224
  signal tmp_ivl_6513 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3225
  signal tmp_ivl_652 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2962
  signal tmp_ivl_6520 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3226
  signal tmp_ivl_6527 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3227
  signal tmp_ivl_653 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2962
  signal tmp_ivl_6534 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3228
  signal tmp_ivl_6536 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3228
  signal tmp_ivl_6543 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3229
  signal tmp_ivl_6545 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3229
  signal tmp_ivl_6552 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3230
  signal tmp_ivl_6554 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3230
  signal tmp_ivl_6561 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3231
  signal tmp_ivl_6563 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3231
  signal tmp_ivl_6570 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3232
  signal tmp_ivl_6572 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3232
  signal tmp_ivl_6579 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3233
  signal tmp_ivl_658 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2962
  signal tmp_ivl_6581 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3233
  signal tmp_ivl_6588 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3234
  signal tmp_ivl_6590 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3234
  signal tmp_ivl_6597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3235
  signal tmp_ivl_6599 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3235
  signal tmp_ivl_660 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2962
  signal tmp_ivl_6606 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3236
  signal tmp_ivl_6608 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3236
  signal tmp_ivl_6615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3237
  signal tmp_ivl_6617 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3237
  signal tmp_ivl_662 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2962
  signal tmp_ivl_6624 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3238
  signal tmp_ivl_6626 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3238
  signal tmp_ivl_6633 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3239
  signal tmp_ivl_6635 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3239
  signal tmp_ivl_6642 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3240
  signal tmp_ivl_6644 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3240
  signal tmp_ivl_6651 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3241
  signal tmp_ivl_6653 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3241
  signal tmp_ivl_6660 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3242
  signal tmp_ivl_6662 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3242
  signal tmp_ivl_6669 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3243
  signal tmp_ivl_6671 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3243
  signal tmp_ivl_6678 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3244
  signal tmp_ivl_668 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2963
  signal tmp_ivl_6680 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3244
  signal tmp_ivl_6687 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3245
  signal tmp_ivl_6689 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3245
  signal tmp_ivl_6696 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3246
  signal tmp_ivl_6698 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3246
  signal tmp_ivl_67 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2942
  signal tmp_ivl_670 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2963
  signal tmp_ivl_6705 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3247
  signal tmp_ivl_6707 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3247
  signal tmp_ivl_671 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2963
  signal tmp_ivl_6714 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3248
  signal tmp_ivl_6716 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3248
  signal tmp_ivl_6723 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3249
  signal tmp_ivl_6725 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3249
  signal tmp_ivl_6732 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3250
  signal tmp_ivl_6734 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3250
  signal tmp_ivl_6741 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3251
  signal tmp_ivl_6743 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3251
  signal tmp_ivl_6750 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3252
  signal tmp_ivl_6752 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3252
  signal tmp_ivl_6759 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3253
  signal tmp_ivl_676 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2963
  signal tmp_ivl_6761 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3253
  signal tmp_ivl_6768 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3254
  signal tmp_ivl_6770 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3254
  signal tmp_ivl_6777 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3255
  signal tmp_ivl_6779 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3255
  signal tmp_ivl_6786 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3256
  signal tmp_ivl_6788 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3256
  signal tmp_ivl_679 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2963
  signal tmp_ivl_6795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3257
  signal tmp_ivl_6797 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3257
  signal tmp_ivl_6804 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3258
  signal tmp_ivl_6806 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3258
  signal tmp_ivl_681 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2963
  signal tmp_ivl_6813 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3259
  signal tmp_ivl_6815 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3259
  signal tmp_ivl_682 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2963
  signal tmp_ivl_6822 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3260
  signal tmp_ivl_6824 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3260
  signal tmp_ivl_6831 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3261
  signal tmp_ivl_6833 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3261
  signal tmp_ivl_6840 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3262
  signal tmp_ivl_6842 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3262
  signal tmp_ivl_6849 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3263
  signal tmp_ivl_6851 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3263
  signal tmp_ivl_6858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3264
  signal tmp_ivl_6860 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3264
  signal tmp_ivl_6867 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3265
  signal tmp_ivl_6869 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3265
  signal tmp_ivl_687 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2963
  signal tmp_ivl_6876 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3266
  signal tmp_ivl_6878 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3266
  signal tmp_ivl_6885 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3267
  signal tmp_ivl_6887 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3267
  signal tmp_ivl_689 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2963
  signal tmp_ivl_6894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3268
  signal tmp_ivl_6896 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3268
  signal tmp_ivl_6903 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3269
  signal tmp_ivl_6905 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3269
  signal tmp_ivl_691 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2963
  signal tmp_ivl_6912 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3270
  signal tmp_ivl_6914 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3270
  signal tmp_ivl_6921 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3271
  signal tmp_ivl_6923 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3271
  signal tmp_ivl_6930 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3272
  signal tmp_ivl_6932 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3272
  signal tmp_ivl_6939 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3273
  signal tmp_ivl_6941 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3273
  signal tmp_ivl_6948 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3274
  signal tmp_ivl_6950 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3274
  signal tmp_ivl_6957 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3275
  signal tmp_ivl_6959 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3275
  signal tmp_ivl_6966 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3276
  signal tmp_ivl_6968 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3276
  signal tmp_ivl_697 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2964
  signal tmp_ivl_6975 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3277
  signal tmp_ivl_6977 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3277
  signal tmp_ivl_6984 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3278
  signal tmp_ivl_6986 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3278
  signal tmp_ivl_699 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2964
  signal tmp_ivl_6993 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3279
  signal tmp_ivl_6995 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3279
  signal tmp_ivl_70 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2942
  signal tmp_ivl_700 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2964
  signal tmp_ivl_7002 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3280
  signal tmp_ivl_7004 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3280
  signal tmp_ivl_7011 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3281
  signal tmp_ivl_7013 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3281
  signal tmp_ivl_7020 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3282
  signal tmp_ivl_7022 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3282
  signal tmp_ivl_7029 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3283
  signal tmp_ivl_7031 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3283
  signal tmp_ivl_7038 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3284
  signal tmp_ivl_7040 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3284
  signal tmp_ivl_7047 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3285
  signal tmp_ivl_7049 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3285
  signal tmp_ivl_705 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2964
  signal tmp_ivl_7056 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3286
  signal tmp_ivl_7058 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3286
  signal tmp_ivl_7065 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3287
  signal tmp_ivl_7067 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3287
  signal tmp_ivl_7074 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3288
  signal tmp_ivl_7076 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3288
  signal tmp_ivl_708 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2964
  signal tmp_ivl_7083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3289
  signal tmp_ivl_7085 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3289
  signal tmp_ivl_7092 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3290
  signal tmp_ivl_7094 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3290
  signal tmp_ivl_710 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2964
  signal tmp_ivl_7101 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3291
  signal tmp_ivl_7103 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3291
  signal tmp_ivl_711 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2964
  signal tmp_ivl_7110 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3292
  signal tmp_ivl_7112 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3292
  signal tmp_ivl_7119 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3293
  signal tmp_ivl_7121 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3293
  signal tmp_ivl_7128 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3294
  signal tmp_ivl_7130 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3294
  signal tmp_ivl_7137 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3295
  signal tmp_ivl_7139 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3295
  signal tmp_ivl_7146 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3296
  signal tmp_ivl_7148 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3296
  signal tmp_ivl_7155 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3297
  signal tmp_ivl_7157 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3297
  signal tmp_ivl_716 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2964
  signal tmp_ivl_7164 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3298
  signal tmp_ivl_7166 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3298
  signal tmp_ivl_7173 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3299
  signal tmp_ivl_7175 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3299
  signal tmp_ivl_718 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2964
  signal tmp_ivl_7182 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3300
  signal tmp_ivl_7184 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3300
  signal tmp_ivl_7191 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3301
  signal tmp_ivl_7193 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3301
  signal tmp_ivl_72 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2942
  signal tmp_ivl_720 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2964
  signal tmp_ivl_7200 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3302
  signal tmp_ivl_7202 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3302
  signal tmp_ivl_7209 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3303
  signal tmp_ivl_7211 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3303
  signal tmp_ivl_7218 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3304
  signal tmp_ivl_7220 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3304
  signal tmp_ivl_7227 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3305
  signal tmp_ivl_7229 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3305
  signal tmp_ivl_7236 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3306
  signal tmp_ivl_7238 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3306
  signal tmp_ivl_7245 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3307
  signal tmp_ivl_7247 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3307
  signal tmp_ivl_7254 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3308
  signal tmp_ivl_7256 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3308
  signal tmp_ivl_726 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2965
  signal tmp_ivl_7263 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3309
  signal tmp_ivl_7265 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3309
  signal tmp_ivl_7272 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3310
  signal tmp_ivl_7274 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3310
  signal tmp_ivl_728 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2965
  signal tmp_ivl_7281 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3311
  signal tmp_ivl_7283 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3311
  signal tmp_ivl_729 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2965
  signal tmp_ivl_7290 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3312
  signal tmp_ivl_7292 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3312
  signal tmp_ivl_7299 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3313
  signal tmp_ivl_73 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2942
  signal tmp_ivl_7301 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3313
  signal tmp_ivl_7308 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3314
  signal tmp_ivl_7310 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3314
  signal tmp_ivl_7317 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3315
  signal tmp_ivl_7319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3315
  signal tmp_ivl_7326 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3316
  signal tmp_ivl_7328 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3316
  signal tmp_ivl_7335 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3317
  signal tmp_ivl_7337 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3317
  signal tmp_ivl_734 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2965
  signal tmp_ivl_7344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3318
  signal tmp_ivl_7346 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3318
  signal tmp_ivl_7353 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3319
  signal tmp_ivl_7355 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3319
  signal tmp_ivl_7362 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3320
  signal tmp_ivl_7364 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3320
  signal tmp_ivl_737 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2965
  signal tmp_ivl_7371 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3321
  signal tmp_ivl_7373 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3321
  signal tmp_ivl_7380 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3322
  signal tmp_ivl_7382 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3322
  signal tmp_ivl_7389 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3323
  signal tmp_ivl_739 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2965
  signal tmp_ivl_7391 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3323
  signal tmp_ivl_7398 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3324
  signal tmp_ivl_740 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2965
  signal tmp_ivl_7400 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3324
  signal tmp_ivl_7407 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3325
  signal tmp_ivl_7409 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3325
  signal tmp_ivl_7416 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3326
  signal tmp_ivl_7418 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3326
  signal tmp_ivl_7425 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3327
  signal tmp_ivl_7427 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3327
  signal tmp_ivl_7434 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3328
  signal tmp_ivl_7436 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3328
  signal tmp_ivl_7443 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3329
  signal tmp_ivl_7445 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3329
  signal tmp_ivl_745 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2965
  signal tmp_ivl_7452 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3330
  signal tmp_ivl_7454 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3330
  signal tmp_ivl_7461 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3331
  signal tmp_ivl_7463 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3331
  signal tmp_ivl_747 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2965
  signal tmp_ivl_7470 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3332
  signal tmp_ivl_7472 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3332
  signal tmp_ivl_7479 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3333
  signal tmp_ivl_7481 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3333
  signal tmp_ivl_7488 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3334
  signal tmp_ivl_749 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2965
  signal tmp_ivl_7490 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3334
  signal tmp_ivl_7497 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3335
  signal tmp_ivl_7499 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3335
  signal tmp_ivl_7506 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3336
  signal tmp_ivl_7508 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3336
  signal tmp_ivl_7515 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3337
  signal tmp_ivl_7517 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3337
  signal tmp_ivl_7524 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3338
  signal tmp_ivl_7526 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3338
  signal tmp_ivl_7533 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3339
  signal tmp_ivl_7535 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3339
  signal tmp_ivl_7542 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3340
  signal tmp_ivl_7544 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3340
  signal tmp_ivl_755 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2966
  signal tmp_ivl_7551 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3341
  signal tmp_ivl_7553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3341
  signal tmp_ivl_7560 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3342
  signal tmp_ivl_7562 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3342
  signal tmp_ivl_7569 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3343
  signal tmp_ivl_757 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2966
  signal tmp_ivl_7571 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3343
  signal tmp_ivl_7578 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3344
  signal tmp_ivl_758 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2966
  signal tmp_ivl_7580 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3344
  signal tmp_ivl_7587 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3345
  signal tmp_ivl_7589 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3345
  signal tmp_ivl_7596 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3346
  signal tmp_ivl_7598 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3346
  signal tmp_ivl_7605 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3347
  signal tmp_ivl_7607 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3347
  signal tmp_ivl_7614 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3348
  signal tmp_ivl_7616 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3348
  signal tmp_ivl_7623 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3349
  signal tmp_ivl_7625 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3349
  signal tmp_ivl_763 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2966
  signal tmp_ivl_7632 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3350
  signal tmp_ivl_7634 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3350
  signal tmp_ivl_7641 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3351
  signal tmp_ivl_7643 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3351
  signal tmp_ivl_7650 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3352
  signal tmp_ivl_7652 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3352
  signal tmp_ivl_7659 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3353
  signal tmp_ivl_766 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2966
  signal tmp_ivl_7661 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3353
  signal tmp_ivl_7668 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3354
  signal tmp_ivl_7670 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3354
  signal tmp_ivl_7677 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3355
  signal tmp_ivl_7679 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3355
  signal tmp_ivl_768 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2966
  signal tmp_ivl_7686 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3361
  signal tmp_ivl_7688 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3361
  signal tmp_ivl_7689 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3361
  signal tmp_ivl_769 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2966
  signal tmp_ivl_7694 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3361
  signal tmp_ivl_7697 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3361
  signal tmp_ivl_7698 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3361
  signal tmp_ivl_7703 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3361
  signal tmp_ivl_7705 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3361
  signal tmp_ivl_7711 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3362
  signal tmp_ivl_7713 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3362
  signal tmp_ivl_7714 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3362
  signal tmp_ivl_7719 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3362
  signal tmp_ivl_7721 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3362
  signal tmp_ivl_7726 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3362
  signal tmp_ivl_7728 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3362
  signal tmp_ivl_7734 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3363
  signal tmp_ivl_7736 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3363
  signal tmp_ivl_7737 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3363
  signal tmp_ivl_774 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2966
  signal tmp_ivl_7742 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3363
  signal tmp_ivl_7745 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3363
  signal tmp_ivl_7746 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3363
  signal tmp_ivl_7751 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3363
  signal tmp_ivl_7753 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3363
  signal tmp_ivl_7759 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3364
  signal tmp_ivl_776 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2966
  signal tmp_ivl_7761 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3364
  signal tmp_ivl_7762 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3364
  signal tmp_ivl_7767 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3364
  signal tmp_ivl_7769 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3364
  signal tmp_ivl_7774 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3364
  signal tmp_ivl_7776 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3364
  signal tmp_ivl_778 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2966
  signal tmp_ivl_7781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3365
  signal tmp_ivl_7786 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3365
  signal tmp_ivl_7788 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3365
  signal tmp_ivl_7793 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3365
  signal tmp_ivl_7795 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3365
  signal tmp_ivl_78 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2942
  signal tmp_ivl_7801 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3366
  signal tmp_ivl_7803 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3366
  signal tmp_ivl_7804 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3366
  signal tmp_ivl_7809 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3366
  signal tmp_ivl_7812 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3366
  signal tmp_ivl_7813 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3366
  signal tmp_ivl_7818 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3366
  signal tmp_ivl_7820 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3366
  signal tmp_ivl_7826 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3367
  signal tmp_ivl_7828 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3367
  signal tmp_ivl_7829 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3367
  signal tmp_ivl_7834 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3367
  signal tmp_ivl_7836 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3367
  signal tmp_ivl_784 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2967
  signal tmp_ivl_7841 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3367
  signal tmp_ivl_7843 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3367
  signal tmp_ivl_7848 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3368
  signal tmp_ivl_7853 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3368
  signal tmp_ivl_7855 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3368
  signal tmp_ivl_786 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2967
  signal tmp_ivl_7860 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3368
  signal tmp_ivl_7862 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3368
  signal tmp_ivl_7864 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3368
  signal tmp_ivl_7866 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3368
  signal tmp_ivl_787 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2967
  signal tmp_ivl_7872 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3369
  signal tmp_ivl_7874 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3369
  signal tmp_ivl_7875 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3369
  signal tmp_ivl_7880 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3369
  signal tmp_ivl_7883 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3369
  signal tmp_ivl_7884 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3369
  signal tmp_ivl_7889 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3369
  signal tmp_ivl_7891 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3369
  signal tmp_ivl_7897 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3370
  signal tmp_ivl_7899 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3370
  signal tmp_ivl_7900 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3370
  signal tmp_ivl_7905 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3370
  signal tmp_ivl_7907 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3370
  signal tmp_ivl_7912 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3370
  signal tmp_ivl_7914 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3370
  signal tmp_ivl_792 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2967
  signal tmp_ivl_7920 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3371
  signal tmp_ivl_7922 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3371
  signal tmp_ivl_7923 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3371
  signal tmp_ivl_7928 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3371
  signal tmp_ivl_7931 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3371
  signal tmp_ivl_7932 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3371
  signal tmp_ivl_7937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3371
  signal tmp_ivl_7939 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3371
  signal tmp_ivl_7945 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3372
  signal tmp_ivl_7947 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3372
  signal tmp_ivl_7948 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3372
  signal tmp_ivl_795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2967
  signal tmp_ivl_7953 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3372
  signal tmp_ivl_7955 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3372
  signal tmp_ivl_7960 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3372
  signal tmp_ivl_7962 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3372
  signal tmp_ivl_7967 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3373
  signal tmp_ivl_797 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2967
  signal tmp_ivl_7972 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3373
  signal tmp_ivl_7974 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3373
  signal tmp_ivl_7979 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3373
  signal tmp_ivl_798 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2967
  signal tmp_ivl_7981 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3373
  signal tmp_ivl_7987 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3374
  signal tmp_ivl_7989 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3374
  signal tmp_ivl_7990 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3374
  signal tmp_ivl_7995 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3374
  signal tmp_ivl_7998 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3374
  signal tmp_ivl_7999 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3374
  signal tmp_ivl_80 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2942
  signal tmp_ivl_8004 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3374
  signal tmp_ivl_8006 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3374
  signal tmp_ivl_8012 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3375
  signal tmp_ivl_8014 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3375
  signal tmp_ivl_8015 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3375
  signal tmp_ivl_8020 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3375
  signal tmp_ivl_8022 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3375
  signal tmp_ivl_8027 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3375
  signal tmp_ivl_8029 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3375
  signal tmp_ivl_803 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2967
  signal tmp_ivl_8034 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3376
  signal tmp_ivl_8039 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3376
  signal tmp_ivl_8041 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3376
  signal tmp_ivl_8046 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3376
  signal tmp_ivl_8048 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3376
  signal tmp_ivl_805 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2967
  signal tmp_ivl_8050 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3376
  signal tmp_ivl_8052 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3376
  signal tmp_ivl_8058 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3377
  signal tmp_ivl_8060 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3377
  signal tmp_ivl_8061 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3377
  signal tmp_ivl_8066 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3377
  signal tmp_ivl_8069 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3377
  signal tmp_ivl_807 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2967
  signal tmp_ivl_8070 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3377
  signal tmp_ivl_8075 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3377
  signal tmp_ivl_8077 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3377
  signal tmp_ivl_8083 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3378
  signal tmp_ivl_8085 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3378
  signal tmp_ivl_8086 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3378
  signal tmp_ivl_8091 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3378
  signal tmp_ivl_8093 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3378
  signal tmp_ivl_8098 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3378
  signal tmp_ivl_8100 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3378
  signal tmp_ivl_8106 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3379
  signal tmp_ivl_8108 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3379
  signal tmp_ivl_8109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3379
  signal tmp_ivl_8114 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3379
  signal tmp_ivl_8117 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3379
  signal tmp_ivl_8118 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3379
  signal tmp_ivl_8123 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3379
  signal tmp_ivl_8125 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3379
  signal tmp_ivl_813 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2968
  signal tmp_ivl_8131 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3380
  signal tmp_ivl_8133 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3380
  signal tmp_ivl_8134 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3380
  signal tmp_ivl_8139 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3380
  signal tmp_ivl_8141 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3380
  signal tmp_ivl_8146 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3380
  signal tmp_ivl_8148 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3380
  signal tmp_ivl_815 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2968
  signal tmp_ivl_8153 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3381
  signal tmp_ivl_8158 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3381
  signal tmp_ivl_816 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2968
  signal tmp_ivl_8160 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3381
  signal tmp_ivl_8165 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3381
  signal tmp_ivl_8167 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3381
  signal tmp_ivl_8173 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3382
  signal tmp_ivl_8175 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3382
  signal tmp_ivl_8176 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3382
  signal tmp_ivl_8181 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3382
  signal tmp_ivl_8184 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3382
  signal tmp_ivl_8185 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3382
  signal tmp_ivl_8190 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3382
  signal tmp_ivl_8192 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3382
  signal tmp_ivl_8198 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3383
  signal tmp_ivl_82 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2942
  signal tmp_ivl_8200 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3383
  signal tmp_ivl_8201 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3383
  signal tmp_ivl_8206 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3383
  signal tmp_ivl_8208 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3383
  signal tmp_ivl_821 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2968
  signal tmp_ivl_8213 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3383
  signal tmp_ivl_8215 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3383
  signal tmp_ivl_8220 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3384
  signal tmp_ivl_8225 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3384
  signal tmp_ivl_8227 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3384
  signal tmp_ivl_8232 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3384
  signal tmp_ivl_8234 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3384
  signal tmp_ivl_8236 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3384
  signal tmp_ivl_8238 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3384
  signal tmp_ivl_824 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2968
  signal tmp_ivl_8244 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3385
  signal tmp_ivl_8246 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3385
  signal tmp_ivl_8247 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3385
  signal tmp_ivl_8252 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3385
  signal tmp_ivl_8255 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3385
  signal tmp_ivl_8256 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3385
  signal tmp_ivl_826 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2968
  signal tmp_ivl_8261 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3385
  signal tmp_ivl_8263 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3385
  signal tmp_ivl_8269 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3386
  signal tmp_ivl_827 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2968
  signal tmp_ivl_8271 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3386
  signal tmp_ivl_8272 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3386
  signal tmp_ivl_8277 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3386
  signal tmp_ivl_8279 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3386
  signal tmp_ivl_8284 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3386
  signal tmp_ivl_8286 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3386
  signal tmp_ivl_8292 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3387
  signal tmp_ivl_8294 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3387
  signal tmp_ivl_8295 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3387
  signal tmp_ivl_8300 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3387
  signal tmp_ivl_8303 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3387
  signal tmp_ivl_8304 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3387
  signal tmp_ivl_8309 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3387
  signal tmp_ivl_8311 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3387
  signal tmp_ivl_8317 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3388
  signal tmp_ivl_8319 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3388
  signal tmp_ivl_832 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2968
  signal tmp_ivl_8320 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3388
  signal tmp_ivl_8325 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3388
  signal tmp_ivl_8327 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3388
  signal tmp_ivl_8332 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3388
  signal tmp_ivl_8334 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3388
  signal tmp_ivl_8339 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3389
  signal tmp_ivl_834 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2968
  signal tmp_ivl_8344 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3389
  signal tmp_ivl_8346 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3389
  signal tmp_ivl_8351 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3389
  signal tmp_ivl_8353 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3389
  signal tmp_ivl_8359 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3390
  signal tmp_ivl_836 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2968
  signal tmp_ivl_8361 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3390
  signal tmp_ivl_8362 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3390
  signal tmp_ivl_8367 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3390
  signal tmp_ivl_8370 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3390
  signal tmp_ivl_8371 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3390
  signal tmp_ivl_8376 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3390
  signal tmp_ivl_8378 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3390
  signal tmp_ivl_8384 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3391
  signal tmp_ivl_8386 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3391
  signal tmp_ivl_8387 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3391
  signal tmp_ivl_8392 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3391
  signal tmp_ivl_8394 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3391
  signal tmp_ivl_8399 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3391
  signal tmp_ivl_8401 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3391
  signal tmp_ivl_8406 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3392
  signal tmp_ivl_8411 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3392
  signal tmp_ivl_8413 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3392
  signal tmp_ivl_8418 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3392
  signal tmp_ivl_842 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2969
  signal tmp_ivl_8420 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3392
  signal tmp_ivl_8422 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3392
  signal tmp_ivl_8424 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3392
  signal tmp_ivl_8430 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3393
  signal tmp_ivl_8432 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3393
  signal tmp_ivl_8433 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3393
  signal tmp_ivl_8438 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3393
  signal tmp_ivl_844 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2969
  signal tmp_ivl_8441 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3393
  signal tmp_ivl_8442 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3393
  signal tmp_ivl_8447 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3393
  signal tmp_ivl_8449 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3393
  signal tmp_ivl_845 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2969
  signal tmp_ivl_8455 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3394
  signal tmp_ivl_8457 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3394
  signal tmp_ivl_8458 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3394
  signal tmp_ivl_8463 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3394
  signal tmp_ivl_8465 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3394
  signal tmp_ivl_8470 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3394
  signal tmp_ivl_8472 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3394
  signal tmp_ivl_8478 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3395
  signal tmp_ivl_8480 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3395
  signal tmp_ivl_8481 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3395
  signal tmp_ivl_8486 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3395
  signal tmp_ivl_8489 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3395
  signal tmp_ivl_8490 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3395
  signal tmp_ivl_8495 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3395
  signal tmp_ivl_8497 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3395
  signal tmp_ivl_850 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2969
  signal tmp_ivl_8503 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3396
  signal tmp_ivl_8505 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3396
  signal tmp_ivl_8506 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3396
  signal tmp_ivl_8511 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3396
  signal tmp_ivl_8513 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3396
  signal tmp_ivl_8518 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3396
  signal tmp_ivl_8520 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3396
  signal tmp_ivl_8525 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3397
  signal tmp_ivl_853 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2969
  signal tmp_ivl_8530 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3397
  signal tmp_ivl_8532 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3397
  signal tmp_ivl_8537 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3397
  signal tmp_ivl_8539 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3397
  signal tmp_ivl_8545 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3398
  signal tmp_ivl_8547 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3398
  signal tmp_ivl_8548 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3398
  signal tmp_ivl_855 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2969
  signal tmp_ivl_8553 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3398
  signal tmp_ivl_8556 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3398
  signal tmp_ivl_8557 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3398
  signal tmp_ivl_856 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2969
  signal tmp_ivl_8562 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3398
  signal tmp_ivl_8564 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3398
  signal tmp_ivl_8570 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3399
  signal tmp_ivl_8572 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3399
  signal tmp_ivl_8573 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3399
  signal tmp_ivl_8578 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3399
  signal tmp_ivl_8580 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3399
  signal tmp_ivl_8585 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3399
  signal tmp_ivl_8587 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3399
  signal tmp_ivl_8592 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3400
  signal tmp_ivl_8597 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3400
  signal tmp_ivl_8599 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3400
  signal tmp_ivl_8604 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3400
  signal tmp_ivl_8606 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3400
  signal tmp_ivl_8608 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3400
  signal tmp_ivl_861 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2969
  signal tmp_ivl_8610 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3400
  signal tmp_ivl_8616 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3401
  signal tmp_ivl_8618 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3401
  signal tmp_ivl_8619 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3401
  signal tmp_ivl_8624 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3401
  signal tmp_ivl_8627 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3401
  signal tmp_ivl_8628 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3401
  signal tmp_ivl_863 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2969
  signal tmp_ivl_8633 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3401
  signal tmp_ivl_8635 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3401
  signal tmp_ivl_8641 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3402
  signal tmp_ivl_8643 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3402
  signal tmp_ivl_8644 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3402
  signal tmp_ivl_8649 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3402
  signal tmp_ivl_865 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2969
  signal tmp_ivl_8651 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3402
  signal tmp_ivl_8656 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3402
  signal tmp_ivl_8658 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3402
  signal tmp_ivl_8664 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3403
  signal tmp_ivl_8666 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3403
  signal tmp_ivl_8667 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3403
  signal tmp_ivl_8672 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3403
  signal tmp_ivl_8675 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3403
  signal tmp_ivl_8676 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3403
  signal tmp_ivl_8681 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3403
  signal tmp_ivl_8683 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3403
  signal tmp_ivl_8689 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3404
  signal tmp_ivl_8691 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3404
  signal tmp_ivl_8692 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3404
  signal tmp_ivl_8697 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3404
  signal tmp_ivl_8699 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3404
  signal tmp_ivl_8704 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3404
  signal tmp_ivl_8706 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3404
  signal tmp_ivl_871 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2970
  signal tmp_ivl_8711 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3405
  signal tmp_ivl_8716 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3405
  signal tmp_ivl_8718 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3405
  signal tmp_ivl_8723 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3405
  signal tmp_ivl_8725 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3405
  signal tmp_ivl_873 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2970
  signal tmp_ivl_8731 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3406
  signal tmp_ivl_8733 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3406
  signal tmp_ivl_8734 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3406
  signal tmp_ivl_8739 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3406
  signal tmp_ivl_874 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2970
  signal tmp_ivl_8742 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3406
  signal tmp_ivl_8743 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3406
  signal tmp_ivl_8748 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3406
  signal tmp_ivl_8750 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3406
  signal tmp_ivl_8756 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3407
  signal tmp_ivl_8758 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3407
  signal tmp_ivl_8759 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3407
  signal tmp_ivl_8764 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3407
  signal tmp_ivl_8766 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3407
  signal tmp_ivl_8771 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3407
  signal tmp_ivl_8773 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3407
  signal tmp_ivl_8778 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3408
  signal tmp_ivl_8783 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3408
  signal tmp_ivl_8785 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3408
  signal tmp_ivl_879 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2970
  signal tmp_ivl_8790 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3408
  signal tmp_ivl_8792 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3408
  signal tmp_ivl_8794 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3408
  signal tmp_ivl_8796 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3408
  signal tmp_ivl_88 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2943
  signal tmp_ivl_8802 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3409
  signal tmp_ivl_8804 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3409
  signal tmp_ivl_8805 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3409
  signal tmp_ivl_8810 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3409
  signal tmp_ivl_8813 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3409
  signal tmp_ivl_8814 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3409
  signal tmp_ivl_8819 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3409
  signal tmp_ivl_882 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2970
  signal tmp_ivl_8821 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3409
  signal tmp_ivl_8827 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3410
  signal tmp_ivl_8829 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3410
  signal tmp_ivl_8830 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3410
  signal tmp_ivl_8835 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3410
  signal tmp_ivl_8837 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3410
  signal tmp_ivl_884 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2970
  signal tmp_ivl_8842 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3410
  signal tmp_ivl_8844 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3410
  signal tmp_ivl_8849 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3411
  signal tmp_ivl_885 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2970
  signal tmp_ivl_8854 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3411
  signal tmp_ivl_8856 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3411
  signal tmp_ivl_8861 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3411
  signal tmp_ivl_8863 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3411
  signal tmp_ivl_8869 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3412
  signal tmp_ivl_8871 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3412
  signal tmp_ivl_8872 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3412
  signal tmp_ivl_8877 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3412
  signal tmp_ivl_8880 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3412
  signal tmp_ivl_8881 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3412
  signal tmp_ivl_8886 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3412
  signal tmp_ivl_8888 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3412
  signal tmp_ivl_8894 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3413
  signal tmp_ivl_8896 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3413
  signal tmp_ivl_8897 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3413
  signal tmp_ivl_890 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2970
  signal tmp_ivl_8902 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3413
  signal tmp_ivl_8904 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3413
  signal tmp_ivl_8909 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3413
  signal tmp_ivl_8911 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3413
  signal tmp_ivl_8916 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3414
  signal tmp_ivl_892 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2970
  signal tmp_ivl_8921 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3414
  signal tmp_ivl_8923 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3414
  signal tmp_ivl_8928 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3414
  signal tmp_ivl_8930 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3414
  signal tmp_ivl_8932 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3414
  signal tmp_ivl_8934 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3414
  signal tmp_ivl_894 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2970
  signal tmp_ivl_8940 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3415
  signal tmp_ivl_8942 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3415
  signal tmp_ivl_8943 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3415
  signal tmp_ivl_8948 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3415
  signal tmp_ivl_8951 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3415
  signal tmp_ivl_8952 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3415
  signal tmp_ivl_8957 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3415
  signal tmp_ivl_8959 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3415
  signal tmp_ivl_8965 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3416
  signal tmp_ivl_8967 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3416
  signal tmp_ivl_8968 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3416
  signal tmp_ivl_8973 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3416
  signal tmp_ivl_8975 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3416
  signal tmp_ivl_8980 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3416
  signal tmp_ivl_8982 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3416
  signal tmp_ivl_8988 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3417
  signal tmp_ivl_8990 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3417
  signal tmp_ivl_8991 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3417
  signal tmp_ivl_8996 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3417
  signal tmp_ivl_8999 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3417
  signal tmp_ivl_9 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2940
  signal tmp_ivl_90 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2943
  signal tmp_ivl_900 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2971
  signal tmp_ivl_9000 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3417
  signal tmp_ivl_9005 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3417
  signal tmp_ivl_9007 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3417
  signal tmp_ivl_9013 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3418
  signal tmp_ivl_9015 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3418
  signal tmp_ivl_9016 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3418
  signal tmp_ivl_902 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2971
  signal tmp_ivl_9021 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3418
  signal tmp_ivl_9023 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3418
  signal tmp_ivl_9028 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3418
  signal tmp_ivl_903 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2971
  signal tmp_ivl_9030 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3418
  signal tmp_ivl_9035 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3419
  signal tmp_ivl_9040 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3419
  signal tmp_ivl_9042 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3419
  signal tmp_ivl_9047 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3419
  signal tmp_ivl_9049 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3419
  signal tmp_ivl_9055 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3420
  signal tmp_ivl_9057 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3420
  signal tmp_ivl_9058 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3420
  signal tmp_ivl_9063 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3420
  signal tmp_ivl_9066 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3420
  signal tmp_ivl_9067 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3420
  signal tmp_ivl_9072 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3420
  signal tmp_ivl_9074 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3420
  signal tmp_ivl_908 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2971
  signal tmp_ivl_9080 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3421
  signal tmp_ivl_9082 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3421
  signal tmp_ivl_9083 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3421
  signal tmp_ivl_9088 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3421
  signal tmp_ivl_9090 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3421
  signal tmp_ivl_9095 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3421
  signal tmp_ivl_9097 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3421
  signal tmp_ivl_91 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2943
  signal tmp_ivl_9102 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3422
  signal tmp_ivl_9107 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3422
  signal tmp_ivl_9109 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3422
  signal tmp_ivl_911 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2971
  signal tmp_ivl_9114 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3422
  signal tmp_ivl_9116 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3422
  signal tmp_ivl_9118 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3422
  signal tmp_ivl_9120 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3422
  signal tmp_ivl_9126 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3423
  signal tmp_ivl_9128 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3423
  signal tmp_ivl_9129 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3423
  signal tmp_ivl_913 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2971
  signal tmp_ivl_9134 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3423
  signal tmp_ivl_9137 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3423
  signal tmp_ivl_9138 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3423
  signal tmp_ivl_914 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2971
  signal tmp_ivl_9143 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3423
  signal tmp_ivl_9145 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3423
  signal tmp_ivl_9151 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3424
  signal tmp_ivl_9153 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3424
  signal tmp_ivl_9154 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3424
  signal tmp_ivl_9159 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3424
  signal tmp_ivl_9161 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3424
  signal tmp_ivl_9166 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3424
  signal tmp_ivl_9168 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3424
  signal tmp_ivl_9173 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3425
  signal tmp_ivl_9178 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3425
  signal tmp_ivl_9180 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3425
  signal tmp_ivl_9185 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3425
  signal tmp_ivl_9187 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3425
  signal tmp_ivl_919 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2971
  signal tmp_ivl_9193 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3426
  signal tmp_ivl_9195 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3426
  signal tmp_ivl_9196 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3426
  signal tmp_ivl_9201 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3426
  signal tmp_ivl_9204 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3426
  signal tmp_ivl_9205 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3426
  signal tmp_ivl_921 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2971
  signal tmp_ivl_9210 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3426
  signal tmp_ivl_9212 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3426
  signal tmp_ivl_9218 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3427
  signal tmp_ivl_9220 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3427
  signal tmp_ivl_9221 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3427
  signal tmp_ivl_9226 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3427
  signal tmp_ivl_9228 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3427
  signal tmp_ivl_923 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2971
  signal tmp_ivl_9233 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3427
  signal tmp_ivl_9235 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3427
  signal tmp_ivl_9240 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3428
  signal tmp_ivl_9245 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3428
  signal tmp_ivl_9247 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3428
  signal tmp_ivl_9252 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3428
  signal tmp_ivl_9254 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3428
  signal tmp_ivl_9256 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3428
  signal tmp_ivl_9258 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3428
  signal tmp_ivl_9264 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3429
  signal tmp_ivl_9266 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3429
  signal tmp_ivl_9267 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3429
  signal tmp_ivl_9272 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3429
  signal tmp_ivl_9275 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3429
  signal tmp_ivl_9276 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3429
  signal tmp_ivl_9281 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3429
  signal tmp_ivl_9283 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3429
  signal tmp_ivl_9289 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3430
  signal tmp_ivl_929 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2972
  signal tmp_ivl_9291 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3430
  signal tmp_ivl_9292 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3430
  signal tmp_ivl_9297 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3430
  signal tmp_ivl_9299 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3430
  signal tmp_ivl_9304 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3430
  signal tmp_ivl_9306 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3430
  signal tmp_ivl_931 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2972
  signal tmp_ivl_9311 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3431
  signal tmp_ivl_9316 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3431
  signal tmp_ivl_9318 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3431
  signal tmp_ivl_932 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2972
  signal tmp_ivl_9323 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3431
  signal tmp_ivl_9325 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3431
  signal tmp_ivl_9331 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3432
  signal tmp_ivl_9333 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3432
  signal tmp_ivl_9334 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3432
  signal tmp_ivl_9339 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3432
  signal tmp_ivl_9342 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3432
  signal tmp_ivl_9343 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3432
  signal tmp_ivl_9348 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3432
  signal tmp_ivl_9350 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3432
  signal tmp_ivl_9356 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3433
  signal tmp_ivl_9358 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3433
  signal tmp_ivl_9359 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3433
  signal tmp_ivl_9364 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3433
  signal tmp_ivl_9366 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3433
  signal tmp_ivl_937 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2972
  signal tmp_ivl_9371 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3433
  signal tmp_ivl_9373 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3433
  signal tmp_ivl_9378 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3434
  signal tmp_ivl_9383 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3434
  signal tmp_ivl_9385 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3434
  signal tmp_ivl_9390 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3434
  signal tmp_ivl_9392 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3434
  signal tmp_ivl_9394 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3434
  signal tmp_ivl_9396 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3434
  signal tmp_ivl_940 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2972
  signal tmp_ivl_9402 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3435
  signal tmp_ivl_9404 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3435
  signal tmp_ivl_9405 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3435
  signal tmp_ivl_9410 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3435
  signal tmp_ivl_9413 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3435
  signal tmp_ivl_9414 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3435
  signal tmp_ivl_9419 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3435
  signal tmp_ivl_942 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2972
  signal tmp_ivl_9421 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3435
  signal tmp_ivl_9427 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3436
  signal tmp_ivl_9429 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3436
  signal tmp_ivl_943 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2972
  signal tmp_ivl_9430 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3436
  signal tmp_ivl_9435 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3436
  signal tmp_ivl_9437 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3436
  signal tmp_ivl_9442 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3436
  signal tmp_ivl_9444 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3436
  signal tmp_ivl_9449 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3437
  signal tmp_ivl_9454 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3437
  signal tmp_ivl_9456 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3437
  signal tmp_ivl_9461 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3437
  signal tmp_ivl_9463 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3437
  signal tmp_ivl_9469 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3438
  signal tmp_ivl_9471 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3438
  signal tmp_ivl_9472 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3438
  signal tmp_ivl_9477 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3438
  signal tmp_ivl_948 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2972
  signal tmp_ivl_9480 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3438
  signal tmp_ivl_9481 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3438
  signal tmp_ivl_9486 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3438
  signal tmp_ivl_9488 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3438
  signal tmp_ivl_9494 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3439
  signal tmp_ivl_9496 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3439
  signal tmp_ivl_9497 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3439
  signal tmp_ivl_950 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2972
  signal tmp_ivl_9502 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3439
  signal tmp_ivl_9504 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3439
  signal tmp_ivl_9509 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3439
  signal tmp_ivl_9511 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3439
  signal tmp_ivl_9516 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3440
  signal tmp_ivl_952 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2972
  signal tmp_ivl_9521 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3440
  signal tmp_ivl_9523 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3440
  signal tmp_ivl_9528 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3440
  signal tmp_ivl_9530 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3440
  signal tmp_ivl_9532 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3440
  signal tmp_ivl_9534 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3440
  signal tmp_ivl_9540 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3441
  signal tmp_ivl_9542 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3441
  signal tmp_ivl_9543 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3441
  signal tmp_ivl_9548 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3441
  signal tmp_ivl_9551 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3441
  signal tmp_ivl_9552 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3441
  signal tmp_ivl_9557 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3441
  signal tmp_ivl_9559 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3441
  signal tmp_ivl_9565 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3442
  signal tmp_ivl_9567 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3442
  signal tmp_ivl_9568 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3442
  signal tmp_ivl_9573 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3442
  signal tmp_ivl_9575 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3442
  signal tmp_ivl_958 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2973
  signal tmp_ivl_9580 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3442
  signal tmp_ivl_9582 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3442
  signal tmp_ivl_9587 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3443
  signal tmp_ivl_9592 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3443
  signal tmp_ivl_9594 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3443
  signal tmp_ivl_9599 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3443
  signal tmp_ivl_96 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2943
  signal tmp_ivl_960 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2973
  signal tmp_ivl_9601 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3443
  signal tmp_ivl_9607 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3444
  signal tmp_ivl_9609 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3444
  signal tmp_ivl_961 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2973
  signal tmp_ivl_9610 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3444
  signal tmp_ivl_9615 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3444
  signal tmp_ivl_9618 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3444
  signal tmp_ivl_9619 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3444
  signal tmp_ivl_9624 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3444
  signal tmp_ivl_9626 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3444
  signal tmp_ivl_9632 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3445
  signal tmp_ivl_9634 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3445
  signal tmp_ivl_9635 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3445
  signal tmp_ivl_9640 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3445
  signal tmp_ivl_9642 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3445
  signal tmp_ivl_9647 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3445
  signal tmp_ivl_9649 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3445
  signal tmp_ivl_9654 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3446
  signal tmp_ivl_9659 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3446
  signal tmp_ivl_966 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2973
  signal tmp_ivl_9661 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3446
  signal tmp_ivl_9666 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3446
  signal tmp_ivl_9668 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3446
  signal tmp_ivl_9670 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3446
  signal tmp_ivl_9672 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3446
  signal tmp_ivl_9677 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3447
  signal tmp_ivl_9682 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3447
  signal tmp_ivl_9684 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3447
  signal tmp_ivl_9689 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3447
  signal tmp_ivl_969 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2973
  signal tmp_ivl_9691 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3447
  signal tmp_ivl_9697 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3448
  signal tmp_ivl_9699 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3448
  signal tmp_ivl_9700 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3448
  signal tmp_ivl_9705 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3448
  signal tmp_ivl_9708 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3448
  signal tmp_ivl_9709 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3448
  signal tmp_ivl_971 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2973
  signal tmp_ivl_9714 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3448
  signal tmp_ivl_9716 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3448
  signal tmp_ivl_972 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2973
  signal tmp_ivl_9722 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3449
  signal tmp_ivl_9724 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3449
  signal tmp_ivl_9725 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3449
  signal tmp_ivl_9730 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3449
  signal tmp_ivl_9732 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3449
  signal tmp_ivl_9737 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3449
  signal tmp_ivl_9739 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3449
  signal tmp_ivl_9744 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3450
  signal tmp_ivl_9749 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3450
  signal tmp_ivl_9751 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3450
  signal tmp_ivl_9756 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3450
  signal tmp_ivl_9758 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3450
  signal tmp_ivl_9760 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3450
  signal tmp_ivl_9762 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3450
  signal tmp_ivl_9767 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3451
  signal tmp_ivl_977 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2973
  signal tmp_ivl_9772 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3451
  signal tmp_ivl_9774 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3451
  signal tmp_ivl_9779 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3451
  signal tmp_ivl_9781 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3451
  signal tmp_ivl_9787 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3452
  signal tmp_ivl_9789 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3452
  signal tmp_ivl_979 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2973
  signal tmp_ivl_9790 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3452
  signal tmp_ivl_9795 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3452
  signal tmp_ivl_9798 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3452
  signal tmp_ivl_9799 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3452
  signal tmp_ivl_9804 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3452
  signal tmp_ivl_9806 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3452
  signal tmp_ivl_981 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2973
  signal tmp_ivl_9812 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3453
  signal tmp_ivl_9814 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3453
  signal tmp_ivl_9815 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3453
  signal tmp_ivl_9820 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3453
  signal tmp_ivl_9822 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3453
  signal tmp_ivl_9827 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3453
  signal tmp_ivl_9829 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3453
  signal tmp_ivl_9834 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3454
  signal tmp_ivl_9839 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3454
  signal tmp_ivl_9841 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3454
  signal tmp_ivl_9846 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3454
  signal tmp_ivl_9848 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3454
  signal tmp_ivl_9850 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3454
  signal tmp_ivl_9852 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3454
  signal tmp_ivl_9858 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3455
  signal tmp_ivl_9860 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3455
  signal tmp_ivl_9861 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3455
  signal tmp_ivl_9866 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3455
  signal tmp_ivl_9869 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3455
  signal tmp_ivl_987 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2974
  signal tmp_ivl_9870 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3455
  signal tmp_ivl_9875 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3455
  signal tmp_ivl_9877 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3455
  signal tmp_ivl_9883 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3456
  signal tmp_ivl_9885 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3456
  signal tmp_ivl_9886 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3456
  signal tmp_ivl_989 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2974
  signal tmp_ivl_9891 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3456
  signal tmp_ivl_9893 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3456
  signal tmp_ivl_9898 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3456
  signal tmp_ivl_99 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2943
  signal tmp_ivl_990 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2974
  signal tmp_ivl_9900 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3456
  signal tmp_ivl_9905 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3457
  signal tmp_ivl_9910 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3457
  signal tmp_ivl_9912 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3457
  signal tmp_ivl_9917 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3457
  signal tmp_ivl_9919 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3457
  signal tmp_ivl_9925 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3458
  signal tmp_ivl_9927 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3458
  signal tmp_ivl_9928 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3458
  signal tmp_ivl_9933 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3458
  signal tmp_ivl_9936 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3458
  signal tmp_ivl_9937 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3458
  signal tmp_ivl_9942 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3458
  signal tmp_ivl_9944 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3458
  signal tmp_ivl_995 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2974
  signal tmp_ivl_9950 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3459
  signal tmp_ivl_9952 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3459
  signal tmp_ivl_9953 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3459
  signal tmp_ivl_9958 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3459
  signal tmp_ivl_9960 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3459
  signal tmp_ivl_9965 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3459
  signal tmp_ivl_9967 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3459
  signal tmp_ivl_9972 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3460
  signal tmp_ivl_9977 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3460
  signal tmp_ivl_9979 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3460
  signal tmp_ivl_998 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2974
  signal tmp_ivl_9984 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3460
  signal tmp_ivl_9986 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3460
  signal tmp_ivl_9988 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3460
  signal tmp_ivl_9990 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3460
  signal tmp_ivl_9996 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3461
  signal tmp_ivl_9998 : std_logic;  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3461
  signal tmp_ivl_9999 : std_logic_vector(1 downto 0);  -- Temporary created at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3461
  signal n3230 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:16
  signal n3231 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:17
  signal n3232 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:18
  signal n3233 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:19
  signal n3234 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:20
  signal n3235 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:21
  signal n3236 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:22
  signal n3237 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:23
  signal n3238 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:24
  signal n3239 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:25
  signal n3240 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:26
  signal n3241 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:27
  signal n3242 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:28
  signal n3243 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:29
  signal n3244 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:30
  signal n3245 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:31
  signal n3246 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:32
  signal n3247 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:33
  signal n3248 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:34
  signal n3249 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:35
  signal n3250 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:36
  signal n3251 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:37
  signal n3252 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:38
  signal n3253 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:39
  signal n3254 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:40
  signal n3255 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:41
  signal n3256 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:42
  signal n3257 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:43
  signal n3258 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:44
  signal n3259 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:45
  signal n3260 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:46
  signal n3261 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:47
  signal n3262 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:48
  signal n3263 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:49
  signal n3264 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:50
  signal n3265 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:51
  signal n3266 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:52
  signal n3267 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:53
  signal n3268 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:54
  signal n3269 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:55
  signal n3270 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:56
  signal n3271 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:57
  signal n3272 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:58
  signal n3273 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:59
  signal n3274 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:60
  signal n3275 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:61
  signal n3276 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:62
  signal n3277 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:63
  signal n3278 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:64
  signal n3279 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:65
  signal n3280 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:66
  signal n3281 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:67
  signal n3282 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:68
  signal n3283 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:69
  signal n3284 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:70
  signal n3285 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:71
  signal n3286 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:72
  signal n3287 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:73
  signal n3288 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:74
  signal n3289 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:75
  signal n3290 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:76
  signal n3291 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:77
  signal n3292 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:78
  signal n3293 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:79
  signal n3294 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:80
  signal n3295 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:81
  signal n3296 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:82
  signal n3297 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:83
  signal n3298 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:84
  signal n3299 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:85
  signal n3300 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:86
  signal n3301 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:87
  signal n3302 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:88
  signal n3303 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:89
  signal n3304 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:90
  signal n3305 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:91
  signal n3306 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:92
  signal n3307 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:93
  signal n3308 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:94
  signal n3309 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:95
  signal n3310 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:96
  signal n3311 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:97
  signal n3312 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:98
  signal n3313 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:99
  signal n3314 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:100
  signal n3315 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:101
  signal n3316 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:102
  signal n3317 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:103
  signal n3318 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:104
  signal n3319 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:105
  signal n3320 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:106
  signal n3321 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:107
  signal n3322 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:108
  signal n3323 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:109
  signal n3324 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:110
  signal n3325 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:111
  signal n3326 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:112
  signal n3327 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:113
  signal n3328 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:114
  signal n3329 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:115
  signal n3330 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:116
  signal n3331 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:117
  signal n3332 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:118
  signal n3333 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:119
  signal n3334 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:120
  signal n3335 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:121
  signal n3336 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:122
  signal n3337 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:123
  signal n3338 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:124
  signal n3339 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:125
  signal n3340 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:126
  signal n3341 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:127
  signal n3342 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:128
  signal n3343 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:129
  signal n3344 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:130
  signal n3345 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:131
  signal n3346 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:132
  signal n3347 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:133
  signal n3348 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:134
  signal n3349 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:135
  signal n3350 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:136
  signal n3351 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:137
  signal n3352 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:138
  signal n3353 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:139
  signal n3354 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:140
  signal n3355 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:141
  signal n3356 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:142
  signal n3357 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:143
  signal n3358 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:144
  signal n3359 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:145
  signal n3360 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:146
  signal n3361 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:147
  signal n3362 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:148
  signal n3363 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:149
  signal n3364 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:150
  signal n3365 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:151
  signal n3366 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:152
  signal n3367 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:153
  signal n3368 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:154
  signal n3369 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:155
  signal n3370 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:156
  signal n3371 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:157
  signal n3372 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:158
  signal n3373 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:159
  signal n3374 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:160
  signal n3375 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:161
  signal n3376 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:162
  signal n3377 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:163
  signal n3378 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:164
  signal n3379 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:165
  signal n3380 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:166
  signal n3381 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:167
  signal n3382 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:168
  signal n3383 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:169
  signal n3384 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:170
  signal n3385 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:171
  signal n3386 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:172
  signal n3387 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:173
  signal n3388 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:174
  signal n3389 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:175
  signal n3390 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:176
  signal n3391 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:177
  signal n3392 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:178
  signal n3393 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:179
  signal n3394 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:180
  signal n3395 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:181
  signal n3396 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:182
  signal n3397 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:183
  signal n3398 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:184
  signal n3399 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:185
  signal n3400 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:186
  signal n3401 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:187
  signal n3402 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:188
  signal n3403 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:189
  signal n3404 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:190
  signal n3405 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:191
  signal n3406 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:192
  signal n3407 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:193
  signal n3408 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:194
  signal n3409 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:195
  signal n3410 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:196
  signal n3411 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:197
  signal n3412 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:198
  signal n3413 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:199
  signal n3414 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:200
  signal n3415 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:201
  signal n3416 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:202
  signal n3417 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:203
  signal n3418 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:204
  signal n3419 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:205
  signal n3420 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:206
  signal n3421 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:207
  signal n3422 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:208
  signal n3423 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:209
  signal n3424 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:210
  signal n3425 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:211
  signal n3426 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:212
  signal n3427 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:213
  signal n3428 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:214
  signal n3429 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:215
  signal n3430 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:216
  signal n3431 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:217
  signal n3432 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:218
  signal n3433 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:219
  signal n3434 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:220
  signal n3435 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:221
  signal n3436 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:222
  signal n3437 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:223
  signal n3438 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:224
  signal n3439 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:225
  signal n3440 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:226
  signal n3441 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:227
  signal n3442 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:228
  signal n3443 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:229
  signal n3444 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:230
  signal n3445 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:231
  signal n3446 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:232
  signal n3447 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:233
  signal n3448 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:234
  signal n3449 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:235
  signal n3450 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:236
  signal n3451 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:237
  signal n3452 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:238
  signal n3453 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:239
  signal n3454 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:240
  signal n3455 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:241
  signal n3456 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:242
  signal n3457 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:243
  signal n3458 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:244
  signal n3459 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:245
  signal n3460 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:246
  signal n3461 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:247
  signal n3462 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:248
  signal n3463 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:249
  signal n3464 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:250
  signal n3465 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:251
  signal n3466 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:252
  signal n3467 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:253
  signal n3468 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:254
  signal n3469 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:255
  signal n3470 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:256
  signal n3471 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:257
  signal n3472 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:258
  signal n3473 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:259
  signal n3474 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:260
  signal n3475 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:261
  signal n3476 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:262
  signal n3477 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:263
  signal n3478 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:264
  signal n3479 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:265
  signal n3480 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:266
  signal n3481 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:267
  signal n3482 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:268
  signal n3483 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:269
  signal n3484 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:270
  signal n3485 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:271
  signal n3486 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:272
  signal n3487 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:273
  signal n3488 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:274
  signal n3489 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:275
  signal n3490 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:276
  signal n3491 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:277
  signal n3492 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:278
  signal n3493 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:279
  signal n3494 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:280
  signal n3495 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:281
  signal n3496 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:282
  signal n3497 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:283
  signal n3498 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:284
  signal n3499 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:285
  signal n3500 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:286
  signal n3501 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:287
  signal n3502 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:288
  signal n3503 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:289
  signal n3504 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:290
  signal n3505 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:291
  signal n3506 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:292
  signal n3507 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:293
  signal n3508 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:294
  signal n3509 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:295
  signal n3510 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:296
  signal n3511 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:297
  signal n3512 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:298
  signal n3513 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:299
  signal n3514 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:300
  signal n3515 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:301
  signal n3516 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:302
  signal n3517 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:303
  signal n3518 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:304
  signal n3519 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:305
  signal n3520 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:306
  signal n3521 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:307
  signal n3522 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:308
  signal n3523 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:309
  signal n3524 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:310
  signal n3525 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:311
  signal n3526 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:312
  signal n3527 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:313
  signal n3528 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:314
  signal n3529 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:315
  signal n3530 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:316
  signal n3531 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:317
  signal n3532 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:318
  signal n3533 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:319
  signal n3534 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:320
  signal n3535 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:321
  signal n3536 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:322
  signal n3537 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:323
  signal n3538 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:324
  signal n3539 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:325
  signal n3540 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:326
  signal n3541 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:327
  signal n3542 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:328
  signal n3543 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:329
  signal n3544 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:330
  signal n3545 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:331
  signal n3546 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:332
  signal n3547 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:333
  signal n3548 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:334
  signal n3549 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:335
  signal n3550 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:336
  signal n3551 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:337
  signal n3552 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:338
  signal n3553 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:339
  signal n3554 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:340
  signal n3555 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:341
  signal n3556 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:342
  signal n3557 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:343
  signal n3558 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:344
  signal n3559 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:345
  signal n3560 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:346
  signal n3561 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:347
  signal n3562 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:348
  signal n3563 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:349
  signal n3564 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:350
  signal n3565 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:351
  signal n3566 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:352
  signal n3567 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:353
  signal n3568 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:354
  signal n3569 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:355
  signal n3570 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:356
  signal n3571 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:357
  signal n3572 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:358
  signal n3573 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:359
  signal n3574 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:360
  signal n3575 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:361
  signal n3576 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:362
  signal n3577 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:363
  signal n3578 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:364
  signal n3579 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:365
  signal n3580 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:366
  signal n3581 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:367
  signal n3582 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:368
  signal n3583 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:369
  signal n3584 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:370
  signal n3585 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:371
  signal n3586 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:372
  signal n3587 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:373
  signal n3588 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:374
  signal n3589 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:375
  signal n3590 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:376
  signal n3591 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:377
  signal n3592 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:378
  signal n3593 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:379
  signal n3594 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:380
  signal n3595 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:381
  signal n3596 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:382
  signal n3597 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:383
  signal n3598 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:384
  signal n3599 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:385
  signal n3600 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:386
  signal n3601 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:387
  signal n3602 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:388
  signal n3603 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:389
  signal n3604 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:390
  signal n3605 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:391
  signal n3606 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:392
  signal n3607 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:393
  signal n3608 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:394
  signal n3609 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:395
  signal n3610 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:396
  signal n3611 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:397
  signal n3612 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:398
  signal n3613 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:399
  signal n3614 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:400
  signal n3615 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:401
  signal n3616 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:402
  signal n3617 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:403
  signal n3618 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:404
  signal n3619 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:405
  signal n3620 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:406
  signal n3621 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:407
  signal n3622 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:408
  signal n3623 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:409
  signal n3624 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:410
  signal n3625 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:411
  signal n3626 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:412
  signal n3627 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:413
  signal n3628 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:414
  signal n3629 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:415
  signal n3630 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:416
  signal n3631 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:417
  signal n3632 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:418
  signal n3633 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:419
  signal n3634 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:420
  signal n3635 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:421
  signal n3636 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:422
  signal n3637 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:423
  signal n3638 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:424
  signal n3639 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:425
  signal n3640 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:426
  signal n3641 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:427
  signal n3642 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:428
  signal n3643 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:429
  signal n3644 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:430
  signal n3645 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:431
  signal n3646 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:432
  signal n3647 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:433
  signal n3648 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:434
  signal n3649 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:435
  signal n3650 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:436
  signal n3651 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:437
  signal n3652 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:438
  signal n3653 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:439
  signal n3654 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:440
  signal n3655 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:441
  signal n3656 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:442
  signal n3657 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:443
  signal n3658 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:444
  signal n3659 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:445
  signal n3660 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:446
  signal n3661 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:447
  signal n3662 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:448
  signal n3663 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:449
  signal n3664 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:450
  signal n3665 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:451
  signal n3666 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:452
  signal n3667 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:453
  signal n3668 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:454
  signal n3669 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:455
  signal n3670 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:456
  signal n3671 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:457
  signal n3672 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:458
  signal n3673 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:459
  signal n3674 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:460
  signal n3675 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:461
  signal n3676 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:462
  signal n3677 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:463
  signal n3678 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:464
  signal n3679 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:465
  signal n3680 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:466
  signal n3681 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:467
  signal n3682 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:468
  signal n3683 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:469
  signal n3684 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:470
  signal n3685 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:471
  signal n3686 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:472
  signal n3687 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:473
  signal n3688 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:474
  signal n3689 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:475
  signal n3690 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:476
  signal n3691 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:477
  signal n3692 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:478
  signal n3693 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:479
  signal n3694 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:480
  signal n3695 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:481
  signal n3696 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:482
  signal n3697 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:483
  signal n3698 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:484
  signal n3699 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:485
  signal n3700 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:486
  signal n3701 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:487
  signal n3702 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:488
  signal n3703 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:489
  signal n3704 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:490
  signal n3705 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:491
  signal n3706 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:492
  signal n3707 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:493
  signal n3708 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:494
  signal n3709 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:495
  signal n3710 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:496
  signal n3711 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:497
  signal n3712 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:498
  signal n3713 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:499
  signal n3714 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:500
  signal n3715 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:501
  signal n3716 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:502
  signal n3717 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:503
  signal n3718 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:504
  signal n3719 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:505
  signal n3720 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:506
  signal n3721 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:507
  signal n3722 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:508
  signal n3723 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:509
  signal n3724 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:510
  signal n3725 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:511
  signal n3726 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:512
  signal n3727 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:513
  signal n3728 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:514
  signal n3729 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:515
  signal n3730 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:516
  signal n3731 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:517
  signal n3732 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:518
  signal n3733 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:519
  signal n3734 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:520
  signal n3735 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:521
  signal n3736 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:522
  signal n3737 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:523
  signal n3738 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:524
  signal n3739 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:525
  signal n3740 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:526
  signal n3741 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:527
  signal n3742 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:528
  signal n3743 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:529
  signal n3744 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:530
  signal n3745 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:531
  signal n3746 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:532
  signal n3747 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:533
  signal n3748 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:534
  signal n3749 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:535
  signal n3750 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:536
  signal n3751 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:537
  signal n3752 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:538
  signal n3753 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:539
  signal n3754 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:540
  signal n3755 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:541
  signal n3756 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:542
  signal n3757 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:543
  signal n3758 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:544
  signal n3759 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:545
  signal n3760 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:546
  signal n3761 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:547
  signal n3762 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:548
  signal n3763 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:549
  signal n3764 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:550
  signal n3765 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:551
  signal n3766 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:552
  signal n3767 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:553
  signal n3768 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:554
  signal n3769 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:555
  signal n3770 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:556
  signal n3771 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:557
  signal n3772 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:558
  signal n3773 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:559
  signal n3774 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:560
  signal n3775 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:561
  signal n3776 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:562
  signal n3777 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:563
  signal n3778 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:564
  signal n3779 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:565
  signal n3780 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:566
  signal n3781 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:567
  signal n3782 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:568
  signal n3783 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:569
  signal n3784 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:570
  signal n3785 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:571
  signal n3786 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:572
  signal n3787 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:573
  signal n3788 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:574
  signal n3789 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:575
  signal n3790 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:576
  signal n3791 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:577
  signal n3792 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:578
  signal n3793 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:579
  signal n3794 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:580
  signal n3795 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:581
  signal n3796 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:582
  signal n3797 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:583
  signal n3798 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:584
  signal n3799 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:585
  signal n3800 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:586
  signal n3801 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:587
  signal n3802 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:588
  signal n3803 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:589
  signal n3804 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:590
  signal n3805 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:591
  signal n3806 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:592
  signal n3807 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:593
  signal n3808 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:594
  signal n3809 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:595
  signal n3810 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:596
  signal n3811 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:597
  signal n3812 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:598
  signal n3813 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:599
  signal n3814 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:600
  signal n3815 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:601
  signal n3816 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:602
  signal n3817 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:603
  signal n3818 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:604
  signal n3819 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:605
  signal n3820 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:606
  signal n3821 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:607
  signal n3822 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:608
  signal n3823 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:609
  signal n3824 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:610
  signal n3825 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:611
  signal n3826 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:612
  signal n3827 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:613
  signal n3828 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:614
  signal n3829 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:615
  signal n3830 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:616
  signal n3831 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:617
  signal n3832 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:618
  signal n3833 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:619
  signal n3834 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:620
  signal n3835 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:621
  signal n3836 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:622
  signal n3837 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:623
  signal n3838 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:624
  signal n3839 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:625
  signal n3840 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:626
  signal n3841 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:627
  signal n3842 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:628
  signal n3843 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:629
  signal n3844 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:630
  signal n3845 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:631
  signal n3846 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:632
  signal n3847 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:633
  signal n3848 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:634
  signal n3849 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:635
  signal n3850 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:636
  signal n3851 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:637
  signal n3852 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:638
  signal n3853 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:639
  signal n3854 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:640
  signal n3855 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:641
  signal n3856 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:642
  signal n3857 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:643
  signal n3858 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:644
  signal n3859 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:645
  signal n3860 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:646
  signal n3861 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:647
  signal n3862 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:648
  signal n3863 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:649
  signal n3864 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:650
  signal n3865 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:651
  signal n3866 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:652
  signal n3867 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:653
  signal n3868 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:654
  signal n3869 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:655
  signal n3870 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:656
  signal n3871 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:657
  signal n3872 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:658
  signal n3873 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:659
  signal n3874 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:660
  signal n3875 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:661
  signal n3876 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:662
  signal n3877 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:663
  signal n3878 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:664
  signal n3879 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:665
  signal n3880 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:666
  signal n3881 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:667
  signal n3882 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:668
  signal n3883 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:669
  signal n3884 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:670
  signal n3885 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:671
  signal n3886 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:672
  signal n3887 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:673
  signal n3888 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:674
  signal n3889 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:675
  signal n3890 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:676
  signal n3891 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:677
  signal n3892 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:678
  signal n3893 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:679
  signal n3894 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:680
  signal n3895 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:681
  signal n3896 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:682
  signal n3897 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:683
  signal n3898 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:684
  signal n3899 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:685
  signal n3900 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:686
  signal n3901 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:687
  signal n3902 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:688
  signal n3903 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:689
  signal n3904 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:690
  signal n3905 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:691
  signal n3906 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:692
  signal n3907 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:693
  signal n3908 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:694
  signal n3909 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:695
  signal n3910 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:696
  signal n3911 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:697
  signal n3912 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:698
  signal n3913 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:699
  signal n3914 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:700
  signal n3915 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:701
  signal n3916 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:702
  signal n3917 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:703
  signal n3918 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:704
  signal n3919 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:705
  signal n3920 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:706
  signal n3921 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:707
  signal n3922 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:708
  signal n3923 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:709
  signal n3924 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:710
  signal n3925 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:711
  signal n3926 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:712
  signal n3927 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:713
  signal n3928 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:714
  signal n3929 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:715
  signal n3930 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:716
  signal n3931 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:717
  signal n3932 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:718
  signal n3933 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:719
  signal n3934 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:720
  signal n3935 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:721
  signal n3936 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:722
  signal n3937 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:723
  signal n3938 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:724
  signal n3939 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:725
  signal n3940 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:726
  signal n3941 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:727
  signal n3942 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:728
  signal n3943 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:729
  signal n3944 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:730
  signal n3945 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:731
  signal n3946 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:732
  signal n3947 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:733
  signal n3948 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:734
  signal n3949 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:735
  signal n3950 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:736
  signal n3951 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:737
  signal n3952 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:738
  signal n3953 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:739
  signal n3954 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:740
  signal n3955 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:741
  signal n3956 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:742
  signal n3957 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:743
  signal n3958 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:744
  signal n3959 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:745
  signal n3960 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:746
  signal n3961 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:747
  signal n3962 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:748
  signal n3963 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:749
  signal n3964 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:750
  signal n3965 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:751
  signal n3966 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:752
  signal n3967 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:753
  signal n3968 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:754
  signal n3969 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:755
  signal n3970 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:756
  signal n3971 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:757
  signal n3972 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:758
  signal n3973 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:759
  signal n3974 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:760
  signal n3975 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:761
  signal n3976 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:762
  signal n3977 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:763
  signal n3978 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:764
  signal n3979 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:765
  signal n3980 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:766
  signal n3981 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:767
  signal n3982 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:768
  signal n3983 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:769
  signal n3984 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:770
  signal n3985 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:771
  signal n3986 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:772
  signal n3987 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:773
  signal n3988 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:774
  signal n3989 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:775
  signal n3990 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:776
  signal n3991 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:777
  signal n3992 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:778
  signal n3993 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:779
  signal n3994 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:780
  signal n3995 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:781
  signal n3996 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:782
  signal n3997 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:783
  signal n3998 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:784
  signal n3999 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:785
  signal n4000 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:786
  signal n4001 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:787
  signal n4002 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:788
  signal n4003 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:789
  signal n4004 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:790
  signal n4005 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:791
  signal n4006 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:792
  signal n4007 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:793
  signal n4008 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:794
  signal n4009 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:795
  signal n4010 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:796
  signal n4011 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:797
  signal n4012 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:798
  signal n4013 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:799
  signal n4014 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:800
  signal n4015 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:801
  signal n4016 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:802
  signal n4017 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:803
  signal n4018 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:804
  signal n4019 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:805
  signal n4020 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:806
  signal n4021 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:807
  signal n4022 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:808
  signal n4023 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:809
  signal n4024 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:810
  signal n4025 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:811
  signal n4026 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:812
  signal n4027 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:813
  signal n4028 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:814
  signal n4029 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:815
  signal n4030 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:816
  signal n4031 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:817
  signal n4032 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:818
  signal n4033 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:819
  signal n4034 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:820
  signal n4035 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:821
  signal n4036 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:822
  signal n4037 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:823
  signal n4038 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:824
  signal n4039 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:825
  signal n4040 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:826
  signal n4041 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:827
  signal n4042 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:828
  signal n4043 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:829
  signal n4044 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:830
  signal n4045 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:831
  signal n4046 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:832
  signal n4047 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:833
  signal n4048 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:834
  signal n4049 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:835
  signal n4050 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:836
  signal n4051 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:837
  signal n4052 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:838
  signal n4053 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:839
  signal n4054 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:840
  signal n4055 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:841
  signal n4056 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:842
  signal n4057 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:843
  signal n4058 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:844
  signal n4059 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:845
  signal n4060 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:846
  signal n4061 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:847
  signal n4062 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:848
  signal n4063 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:849
  signal n4064 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:850
  signal n4065 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:851
  signal n4066 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:852
  signal n4067 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:853
  signal n4068 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:854
  signal n4069 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:855
  signal n4070 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:856
  signal n4071 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:857
  signal n4072 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:858
  signal n4073 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:859
  signal n4074 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:860
  signal n4075 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:861
  signal n4076 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:862
  signal n4077 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:863
  signal n4078 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:864
  signal n4079 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:865
  signal n4080 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:866
  signal n4081 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:867
  signal n4082 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:868
  signal n4083 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:869
  signal n4084 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:870
  signal n4085 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:871
  signal n4086 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:872
  signal n4087 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:873
  signal n4088 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:874
  signal n4089 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:875
  signal n4090 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:876
  signal n4091 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:877
  signal n4092 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:878
  signal n4093 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:879
  signal n4094 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:880
  signal n4095 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:881
  signal n4096 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:882
  signal n4097 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:883
  signal n4098 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:884
  signal n4099 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:885
  signal n4100 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:886
  signal n4101 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:887
  signal n4102 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:888
  signal n4103 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:889
  signal n4104 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:890
  signal n4105 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:891
  signal n4106 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:892
  signal n4107 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:893
  signal n4108 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:894
  signal n4109 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:895
  signal n4110 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:896
  signal n4111 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:897
  signal n4112 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:898
  signal n4113 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:899
  signal n4114 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:900
  signal n4115 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:901
  signal n4116 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:902
  signal n4117 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:903
  signal n4118 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:904
  signal n4119 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:905
  signal n4120 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:906
  signal n4121 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:907
  signal n4122 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:908
  signal n4123 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:909
  signal n4124 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:910
  signal n4125 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:911
  signal n4126 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:912
  signal n4127 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:913
  signal n4128 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:914
  signal n4129 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:915
  signal n4130 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:916
  signal n4131 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:917
  signal n4132 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:918
  signal n4133 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:919
  signal n4134 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:920
  signal n4135 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:921
  signal n4136 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:922
  signal n4137 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:923
  signal n4138 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:924
  signal n4139 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:925
  signal n4140 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:926
  signal n4141 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:927
  signal n4142 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:928
  signal n4143 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:929
  signal n4144 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:930
  signal n4145 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:931
  signal n4146 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:932
  signal n4147 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:933
  signal n4148 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:934
  signal n4149 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:935
  signal n4150 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:936
  signal n4151 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:937
  signal n4152 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:938
  signal n4153 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:939
  signal n4154 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:940
  signal n4155 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:941
  signal n4156 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:942
  signal n4157 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:943
  signal n4158 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:944
  signal n4159 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:945
  signal n4160 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:946
  signal n4161 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:947
  signal n4162 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:948
  signal n4163 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:949
  signal n4164 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:950
  signal n4165 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:951
  signal n4166 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:952
  signal n4167 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:953
  signal n4168 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:954
  signal n4169 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:955
  signal n4170 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:956
  signal n4171 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:957
  signal n4172 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:958
  signal n4173 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:959
  signal n4174 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:960
  signal n4175 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:961
  signal n4176 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:962
  signal n4177 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:963
  signal n4178 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:964
  signal n4179 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:965
  signal n4180 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:966
  signal n4181 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:967
  signal n4182 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:968
  signal n4183 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:969
  signal n4184 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:970
  signal n4185 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:971
  signal n4186 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:972
  signal n4187 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:973
  signal n4188 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:974
  signal n4189 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:975
  signal n4190 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:976
  signal n4191 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:977
  signal n4192 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:978
  signal n4193 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:979
  signal n4194 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:980
  signal n4195 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:981
  signal n4196 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:982
  signal n4197 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:983
  signal n4198 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:984
  signal n4199 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:985
  signal n4200 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:986
  signal n4201 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:987
  signal n4202 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:988
  signal n4203 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:989
  signal n4204 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:990
  signal n4205 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:991
  signal n4206 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:992
  signal n4207 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:993
  signal n4208 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:994
  signal n4209 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:995
  signal n4210 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:996
  signal n4211 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:997
  signal n4212 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:998
  signal n4213 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:999
  signal n4214 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1000
  signal n4215 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1001
  signal n4216 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1002
  signal n4217 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1003
  signal n4218 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1004
  signal n4219 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1005
  signal n4220 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1006
  signal n4221 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1007
  signal n4222 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1008
  signal n4223 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1009
  signal n4224 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1010
  signal n4225 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1011
  signal n4226 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1012
  signal n4227 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1013
  signal n4228 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1014
  signal n4229 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1015
  signal n4230 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1016
  signal n4231 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1017
  signal n4232 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1018
  signal n4233 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1019
  signal n4234 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1020
  signal n4235 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1021
  signal n4236 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1022
  signal n4237 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1023
  signal n4238 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1024
  signal n4239 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1025
  signal n4240 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1026
  signal n4241 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1027
  signal n4242 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1028
  signal n4243 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1029
  signal n4244 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1030
  signal n4245 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1031
  signal n4246 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1032
  signal n4247 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1033
  signal n4248 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1034
  signal n4249 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1035
  signal n4250 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1036
  signal n4251 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1037
  signal n4252 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1038
  signal n4253 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1039
  signal n4254 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1040
  signal n4255 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1041
  signal n4256 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1042
  signal n4257 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1043
  signal n4258 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1044
  signal n4259 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1045
  signal n4260 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1046
  signal n4261 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1047
  signal n4262 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1048
  signal n4263 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1049
  signal n4264 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1050
  signal n4265 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1051
  signal n4266 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1052
  signal n4267 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1053
  signal n4268 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1054
  signal n4269 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1055
  signal n4270 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1056
  signal n4271 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1057
  signal n4272 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1058
  signal new_AGEMA_signal_2338 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1259
  signal new_AGEMA_signal_2341 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1260
  signal new_AGEMA_signal_2344 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1261
  signal new_AGEMA_signal_2347 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1262
  signal new_AGEMA_signal_2350 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1263
  signal new_AGEMA_signal_2353 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1264
  signal new_AGEMA_signal_2356 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1265
  signal new_AGEMA_signal_2359 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1266
  signal new_AGEMA_signal_2362 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1267
  signal new_AGEMA_signal_2365 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1268
  signal new_AGEMA_signal_2368 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1269
  signal new_AGEMA_signal_2371 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1270
  signal new_AGEMA_signal_2374 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1271
  signal new_AGEMA_signal_2377 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1272
  signal new_AGEMA_signal_2380 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1273
  signal new_AGEMA_signal_2383 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1274
  signal new_AGEMA_signal_2386 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1275
  signal new_AGEMA_signal_2389 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1276
  signal new_AGEMA_signal_2392 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1277
  signal new_AGEMA_signal_2395 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1278
  signal new_AGEMA_signal_2398 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1279
  signal new_AGEMA_signal_2401 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1280
  signal new_AGEMA_signal_2404 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1281
  signal new_AGEMA_signal_2407 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1282
  signal new_AGEMA_signal_2410 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1283
  signal new_AGEMA_signal_2413 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1284
  signal new_AGEMA_signal_2416 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1285
  signal new_AGEMA_signal_2419 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1286
  signal new_AGEMA_signal_2422 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1287
  signal new_AGEMA_signal_2425 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1288
  signal new_AGEMA_signal_2428 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1289
  signal new_AGEMA_signal_2431 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1290
  signal new_AGEMA_signal_2434 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1291
  signal new_AGEMA_signal_2437 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1292
  signal new_AGEMA_signal_2440 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1293
  signal new_AGEMA_signal_2443 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1294
  signal new_AGEMA_signal_2446 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1295
  signal new_AGEMA_signal_2449 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1296
  signal new_AGEMA_signal_2452 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1297
  signal new_AGEMA_signal_2455 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1298
  signal new_AGEMA_signal_2458 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1299
  signal new_AGEMA_signal_2461 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1300
  signal new_AGEMA_signal_2464 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1301
  signal new_AGEMA_signal_2467 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1302
  signal new_AGEMA_signal_2470 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1303
  signal new_AGEMA_signal_2473 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1304
  signal new_AGEMA_signal_2476 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1305
  signal new_AGEMA_signal_2479 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1306
  signal new_AGEMA_signal_2482 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1307
  signal new_AGEMA_signal_2485 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1308
  signal new_AGEMA_signal_2488 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1309
  signal new_AGEMA_signal_2491 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1310
  signal new_AGEMA_signal_2494 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1311
  signal new_AGEMA_signal_2497 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1312
  signal new_AGEMA_signal_2500 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1313
  signal new_AGEMA_signal_2503 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1314
  signal new_AGEMA_signal_2506 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1315
  signal new_AGEMA_signal_2509 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1316
  signal new_AGEMA_signal_2512 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1317
  signal new_AGEMA_signal_2515 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1318
  signal new_AGEMA_signal_2518 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1319
  signal new_AGEMA_signal_2521 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1320
  signal new_AGEMA_signal_2524 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1321
  signal new_AGEMA_signal_2527 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1322
  signal new_AGEMA_signal_2529 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1323
  signal new_AGEMA_signal_2531 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1324
  signal new_AGEMA_signal_2533 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1325
  signal new_AGEMA_signal_2535 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1326
  signal new_AGEMA_signal_2537 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1327
  signal new_AGEMA_signal_2539 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1328
  signal new_AGEMA_signal_2541 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1329
  signal new_AGEMA_signal_2543 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1330
  signal new_AGEMA_signal_2545 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1331
  signal new_AGEMA_signal_2547 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1332
  signal new_AGEMA_signal_2549 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1333
  signal new_AGEMA_signal_2551 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1334
  signal new_AGEMA_signal_2553 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1335
  signal new_AGEMA_signal_2555 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1336
  signal new_AGEMA_signal_2557 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1337
  signal new_AGEMA_signal_2559 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1338
  signal new_AGEMA_signal_2561 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1339
  signal new_AGEMA_signal_2563 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1340
  signal new_AGEMA_signal_2565 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1341
  signal new_AGEMA_signal_2567 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1342
  signal new_AGEMA_signal_2569 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1343
  signal new_AGEMA_signal_2571 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1344
  signal new_AGEMA_signal_2573 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1345
  signal new_AGEMA_signal_2575 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1346
  signal new_AGEMA_signal_2577 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1347
  signal new_AGEMA_signal_2579 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1348
  signal new_AGEMA_signal_2581 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1349
  signal new_AGEMA_signal_2583 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1350
  signal new_AGEMA_signal_2585 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1351
  signal new_AGEMA_signal_2587 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1352
  signal new_AGEMA_signal_2589 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1353
  signal new_AGEMA_signal_2591 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1354
  signal new_AGEMA_signal_2593 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1355
  signal new_AGEMA_signal_2595 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1356
  signal new_AGEMA_signal_2597 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1357
  signal new_AGEMA_signal_2599 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1358
  signal new_AGEMA_signal_2601 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1359
  signal new_AGEMA_signal_2603 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1360
  signal new_AGEMA_signal_2605 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1361
  signal new_AGEMA_signal_2607 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1362
  signal new_AGEMA_signal_2609 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1363
  signal new_AGEMA_signal_2611 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1364
  signal new_AGEMA_signal_2613 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1365
  signal new_AGEMA_signal_2615 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1366
  signal new_AGEMA_signal_2617 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1367
  signal new_AGEMA_signal_2619 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1368
  signal new_AGEMA_signal_2621 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1369
  signal new_AGEMA_signal_2623 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1370
  signal new_AGEMA_signal_2625 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1371
  signal new_AGEMA_signal_2627 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1372
  signal new_AGEMA_signal_2629 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1373
  signal new_AGEMA_signal_2631 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1374
  signal new_AGEMA_signal_2633 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1375
  signal new_AGEMA_signal_2635 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1376
  signal new_AGEMA_signal_2637 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1377
  signal new_AGEMA_signal_2639 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1378
  signal new_AGEMA_signal_2641 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1379
  signal new_AGEMA_signal_2643 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1380
  signal new_AGEMA_signal_2645 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1381
  signal new_AGEMA_signal_2647 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1382
  signal new_AGEMA_signal_2649 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1383
  signal new_AGEMA_signal_2651 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1384
  signal new_AGEMA_signal_2653 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1385
  signal new_AGEMA_signal_2655 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1386
  signal new_AGEMA_signal_2657 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1387
  signal new_AGEMA_signal_2659 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1388
  signal new_AGEMA_signal_2661 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1389
  signal new_AGEMA_signal_2663 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1390
  signal new_AGEMA_signal_2665 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1391
  signal new_AGEMA_signal_2667 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1392
  signal new_AGEMA_signal_2669 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1393
  signal new_AGEMA_signal_2671 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1394
  signal new_AGEMA_signal_2673 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1395
  signal new_AGEMA_signal_2675 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1396
  signal new_AGEMA_signal_2677 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1397
  signal new_AGEMA_signal_2679 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1398
  signal new_AGEMA_signal_2681 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1399
  signal new_AGEMA_signal_2683 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1400
  signal new_AGEMA_signal_2685 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1401
  signal new_AGEMA_signal_2687 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1402
  signal new_AGEMA_signal_2689 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1403
  signal new_AGEMA_signal_2692 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1404
  signal new_AGEMA_signal_2695 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1405
  signal new_AGEMA_signal_2698 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1406
  signal new_AGEMA_signal_2701 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1407
  signal new_AGEMA_signal_2704 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1408
  signal new_AGEMA_signal_2707 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1409
  signal new_AGEMA_signal_2709 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1410
  signal new_AGEMA_signal_2712 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1411
  signal new_AGEMA_signal_2714 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1412
  signal new_AGEMA_signal_2717 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1413
  signal new_AGEMA_signal_2719 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1414
  signal new_AGEMA_signal_2721 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1415
  signal new_AGEMA_signal_2724 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1416
  signal new_AGEMA_signal_2727 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1417
  signal new_AGEMA_signal_2730 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1418
  signal new_AGEMA_signal_2733 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1419
  signal new_AGEMA_signal_2736 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1420
  signal new_AGEMA_signal_2739 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1421
  signal new_AGEMA_signal_2742 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1422
  signal new_AGEMA_signal_2744 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1423
  signal new_AGEMA_signal_2747 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1424
  signal new_AGEMA_signal_2750 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1425
  signal new_AGEMA_signal_2753 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1426
  signal new_AGEMA_signal_2755 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1427
  signal new_AGEMA_signal_2758 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1428
  signal new_AGEMA_signal_2760 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1429
  signal new_AGEMA_signal_2763 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1430
  signal new_AGEMA_signal_2766 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1431
  signal new_AGEMA_signal_2769 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1432
  signal new_AGEMA_signal_2772 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1433
  signal new_AGEMA_signal_2775 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1434
  signal new_AGEMA_signal_2778 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1435
  signal new_AGEMA_signal_2780 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1436
  signal new_AGEMA_signal_2783 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1437
  signal new_AGEMA_signal_2786 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1438
  signal new_AGEMA_signal_2788 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1439
  signal new_AGEMA_signal_2790 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1440
  signal new_AGEMA_signal_2793 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1441
  signal new_AGEMA_signal_2795 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1442
  signal new_AGEMA_signal_2797 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1443
  signal new_AGEMA_signal_2800 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1444
  signal new_AGEMA_signal_2803 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1445
  signal new_AGEMA_signal_2805 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1446
  signal new_AGEMA_signal_2807 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1447
  signal new_AGEMA_signal_2810 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1448
  signal new_AGEMA_signal_2813 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1449
  signal new_AGEMA_signal_2816 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1450
  signal new_AGEMA_signal_2819 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1451
  signal new_AGEMA_signal_2821 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1452
  signal new_AGEMA_signal_2823 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1453
  signal new_AGEMA_signal_2825 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1454
  signal new_AGEMA_signal_2828 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1455
  signal new_AGEMA_signal_2831 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1456
  signal new_AGEMA_signal_2834 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1457
  signal new_AGEMA_signal_2837 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1458
  signal new_AGEMA_signal_2840 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1459
  signal new_AGEMA_signal_2843 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1460
  signal new_AGEMA_signal_2846 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1461
  signal new_AGEMA_signal_2849 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1462
  signal new_AGEMA_signal_2852 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1463
  signal new_AGEMA_signal_2855 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1464
  signal new_AGEMA_signal_2858 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1465
  signal new_AGEMA_signal_2859 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1466
  signal new_AGEMA_signal_2860 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1467
  signal new_AGEMA_signal_2861 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1468
  signal new_AGEMA_signal_2862 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1469
  signal new_AGEMA_signal_2863 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1470
  signal new_AGEMA_signal_2864 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1471
  signal new_AGEMA_signal_2865 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1472
  signal new_AGEMA_signal_2866 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1473
  signal new_AGEMA_signal_2867 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1474
  signal new_AGEMA_signal_2868 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1475
  signal new_AGEMA_signal_2869 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1476
  signal new_AGEMA_signal_2870 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1477
  signal new_AGEMA_signal_2871 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1478
  signal new_AGEMA_signal_2872 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1479
  signal new_AGEMA_signal_2873 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1480
  signal new_AGEMA_signal_2874 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1481
  signal new_AGEMA_signal_2875 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1482
  signal new_AGEMA_signal_2876 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1483
  signal new_AGEMA_signal_2877 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1484
  signal new_AGEMA_signal_2878 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1485
  signal new_AGEMA_signal_2879 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1486
  signal new_AGEMA_signal_2880 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1487
  signal new_AGEMA_signal_2881 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1488
  signal new_AGEMA_signal_2882 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1489
  signal new_AGEMA_signal_2883 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1490
  signal new_AGEMA_signal_2884 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1491
  signal new_AGEMA_signal_2885 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1492
  signal new_AGEMA_signal_2886 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1493
  signal new_AGEMA_signal_2887 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1494
  signal new_AGEMA_signal_2888 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1495
  signal new_AGEMA_signal_2889 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1496
  signal new_AGEMA_signal_2890 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1497
  signal new_AGEMA_signal_2891 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1498
  signal new_AGEMA_signal_2892 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1499
  signal new_AGEMA_signal_2893 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1500
  signal new_AGEMA_signal_2894 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1501
  signal new_AGEMA_signal_2895 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1502
  signal new_AGEMA_signal_2896 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1503
  signal new_AGEMA_signal_2897 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1504
  signal new_AGEMA_signal_2899 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1505
  signal new_AGEMA_signal_2900 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1506
  signal new_AGEMA_signal_2901 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1507
  signal new_AGEMA_signal_2902 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1508
  signal new_AGEMA_signal_2904 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1509
  signal new_AGEMA_signal_2905 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1510
  signal new_AGEMA_signal_2906 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1511
  signal new_AGEMA_signal_2907 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1512
  signal new_AGEMA_signal_2908 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1513
  signal new_AGEMA_signal_2909 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1514
  signal new_AGEMA_signal_2910 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1515
  signal new_AGEMA_signal_2911 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1516
  signal new_AGEMA_signal_2912 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1517
  signal new_AGEMA_signal_2913 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1518
  signal new_AGEMA_signal_2914 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1519
  signal new_AGEMA_signal_2915 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1520
  signal new_AGEMA_signal_2916 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1521
  signal new_AGEMA_signal_2917 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1522
  signal new_AGEMA_signal_2918 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1523
  signal new_AGEMA_signal_2919 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1524
  signal new_AGEMA_signal_2920 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1525
  signal new_AGEMA_signal_2921 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1526
  signal new_AGEMA_signal_2922 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1527
  signal new_AGEMA_signal_2923 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1528
  signal new_AGEMA_signal_2924 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1529
  signal new_AGEMA_signal_2925 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1530
  signal new_AGEMA_signal_2926 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1531
  signal new_AGEMA_signal_2927 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1532
  signal new_AGEMA_signal_2928 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1533
  signal new_AGEMA_signal_2929 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1534
  signal new_AGEMA_signal_2930 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1535
  signal new_AGEMA_signal_2931 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1536
  signal new_AGEMA_signal_2932 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1537
  signal new_AGEMA_signal_2933 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1538
  signal new_AGEMA_signal_2934 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1539
  signal new_AGEMA_signal_2935 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1540
  signal new_AGEMA_signal_2936 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1541
  signal new_AGEMA_signal_2937 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1542
  signal new_AGEMA_signal_2938 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1543
  signal new_AGEMA_signal_2939 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1544
  signal new_AGEMA_signal_2940 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1545
  signal new_AGEMA_signal_2941 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1546
  signal new_AGEMA_signal_2942 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1547
  signal new_AGEMA_signal_2943 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1548
  signal new_AGEMA_signal_2944 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1549
  signal new_AGEMA_signal_2945 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1550
  signal new_AGEMA_signal_2946 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1551
  signal new_AGEMA_signal_2947 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1552
  signal new_AGEMA_signal_2948 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1553
  signal new_AGEMA_signal_2949 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1554
  signal new_AGEMA_signal_2950 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1555
  signal new_AGEMA_signal_2951 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1556
  signal new_AGEMA_signal_2952 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1557
  signal new_AGEMA_signal_2953 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1558
  signal new_AGEMA_signal_2954 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1559
  signal new_AGEMA_signal_2955 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1560
  signal new_AGEMA_signal_2956 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1561
  signal new_AGEMA_signal_2957 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1562
  signal new_AGEMA_signal_2958 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1563
  signal new_AGEMA_signal_2959 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1564
  signal new_AGEMA_signal_2960 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1565
  signal new_AGEMA_signal_2961 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1566
  signal new_AGEMA_signal_2962 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1567
  signal new_AGEMA_signal_2963 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1568
  signal new_AGEMA_signal_2964 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1569
  signal new_AGEMA_signal_2965 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1570
  signal new_AGEMA_signal_2966 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1571
  signal new_AGEMA_signal_2967 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1572
  signal new_AGEMA_signal_2968 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1573
  signal new_AGEMA_signal_2969 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1574
  signal new_AGEMA_signal_2970 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1575
  signal new_AGEMA_signal_2971 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1576
  signal new_AGEMA_signal_2972 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1577
  signal new_AGEMA_signal_2973 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1578
  signal new_AGEMA_signal_2974 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1579
  signal new_AGEMA_signal_2975 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1580
  signal new_AGEMA_signal_2976 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1581
  signal new_AGEMA_signal_2977 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1582
  signal new_AGEMA_signal_2978 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1583
  signal new_AGEMA_signal_2979 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1584
  signal new_AGEMA_signal_2980 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1585
  signal new_AGEMA_signal_2981 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1586
  signal new_AGEMA_signal_2982 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1587
  signal new_AGEMA_signal_2983 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1588
  signal new_AGEMA_signal_2984 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1589
  signal new_AGEMA_signal_2985 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1590
  signal new_AGEMA_signal_2986 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1591
  signal new_AGEMA_signal_2987 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1592
  signal new_AGEMA_signal_2988 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1593
  signal new_AGEMA_signal_2989 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1594
  signal new_AGEMA_signal_2990 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1595
  signal new_AGEMA_signal_2991 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1596
  signal new_AGEMA_signal_2992 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1597
  signal new_AGEMA_signal_2993 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1598
  signal new_AGEMA_signal_2994 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1599
  signal new_AGEMA_signal_2995 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1600
  signal new_AGEMA_signal_2996 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1601
  signal new_AGEMA_signal_2997 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1602
  signal new_AGEMA_signal_2998 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1603
  signal new_AGEMA_signal_2999 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1604
  signal new_AGEMA_signal_3000 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1605
  signal new_AGEMA_signal_3001 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1606
  signal new_AGEMA_signal_3002 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1607
  signal new_AGEMA_signal_3003 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1608
  signal new_AGEMA_signal_3004 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1609
  signal new_AGEMA_signal_3005 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1610
  signal new_AGEMA_signal_3006 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1611
  signal new_AGEMA_signal_3007 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1612
  signal new_AGEMA_signal_3008 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1613
  signal new_AGEMA_signal_3009 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1614
  signal new_AGEMA_signal_3010 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1615
  signal new_AGEMA_signal_3011 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1616
  signal new_AGEMA_signal_3012 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1617
  signal new_AGEMA_signal_3013 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1618
  signal new_AGEMA_signal_3014 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1619
  signal new_AGEMA_signal_3015 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1620
  signal new_AGEMA_signal_3016 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1621
  signal new_AGEMA_signal_3017 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1622
  signal new_AGEMA_signal_3018 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1623
  signal new_AGEMA_signal_3019 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1624
  signal new_AGEMA_signal_3020 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1625
  signal new_AGEMA_signal_3021 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1626
  signal new_AGEMA_signal_3022 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1627
  signal new_AGEMA_signal_3023 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1628
  signal new_AGEMA_signal_3024 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1629
  signal new_AGEMA_signal_3025 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1630
  signal new_AGEMA_signal_3026 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1631
  signal new_AGEMA_signal_3027 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1632
  signal new_AGEMA_signal_3028 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1633
  signal new_AGEMA_signal_3029 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1634
  signal new_AGEMA_signal_3030 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1635
  signal new_AGEMA_signal_3031 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1636
  signal new_AGEMA_signal_3032 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1637
  signal new_AGEMA_signal_3033 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1638
  signal new_AGEMA_signal_3034 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1639
  signal new_AGEMA_signal_3035 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1640
  signal new_AGEMA_signal_3036 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1641
  signal new_AGEMA_signal_3037 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1642
  signal new_AGEMA_signal_3038 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1643
  signal new_AGEMA_signal_3039 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1644
  signal new_AGEMA_signal_3040 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1645
  signal new_AGEMA_signal_3041 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1646
  signal new_AGEMA_signal_3042 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1647
  signal new_AGEMA_signal_3043 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1648
  signal new_AGEMA_signal_3044 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1649
  signal new_AGEMA_signal_3045 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1650
  signal new_AGEMA_signal_3046 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1651
  signal new_AGEMA_signal_3047 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1652
  signal new_AGEMA_signal_3048 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1653
  signal new_AGEMA_signal_3049 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1654
  signal new_AGEMA_signal_3050 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1655
  signal new_AGEMA_signal_3051 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1656
  signal new_AGEMA_signal_3052 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1657
  signal new_AGEMA_signal_3053 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1658
  signal new_AGEMA_signal_3054 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1659
  signal new_AGEMA_signal_3055 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1660
  signal new_AGEMA_signal_3056 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1661
  signal new_AGEMA_signal_3057 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1662
  signal new_AGEMA_signal_3058 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1663
  signal new_AGEMA_signal_3059 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1664
  signal new_AGEMA_signal_3060 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1665
  signal new_AGEMA_signal_3061 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1666
  signal new_AGEMA_signal_3062 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1667
  signal new_AGEMA_signal_3063 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1668
  signal new_AGEMA_signal_3064 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1669
  signal new_AGEMA_signal_3065 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1670
  signal new_AGEMA_signal_3066 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1671
  signal new_AGEMA_signal_3067 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1672
  signal new_AGEMA_signal_3068 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1673
  signal new_AGEMA_signal_3069 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1674
  signal new_AGEMA_signal_3070 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1675
  signal new_AGEMA_signal_3071 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1676
  signal new_AGEMA_signal_3072 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1677
  signal new_AGEMA_signal_3073 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1678
  signal new_AGEMA_signal_3074 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1679
  signal new_AGEMA_signal_3075 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1680
  signal new_AGEMA_signal_3076 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1681
  signal new_AGEMA_signal_3077 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1682
  signal new_AGEMA_signal_3078 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1683
  signal new_AGEMA_signal_3079 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1684
  signal new_AGEMA_signal_3080 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1685
  signal new_AGEMA_signal_3081 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1686
  signal new_AGEMA_signal_3082 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1687
  signal new_AGEMA_signal_3083 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1688
  signal new_AGEMA_signal_3084 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1689
  signal new_AGEMA_signal_3085 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1690
  signal new_AGEMA_signal_3086 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1691
  signal new_AGEMA_signal_3087 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1692
  signal new_AGEMA_signal_3088 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1693
  signal new_AGEMA_signal_3089 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1694
  signal new_AGEMA_signal_3090 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1695
  signal new_AGEMA_signal_3091 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1696
  signal new_AGEMA_signal_3092 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1697
  signal new_AGEMA_signal_3093 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1698
  signal new_AGEMA_signal_3094 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1699
  signal new_AGEMA_signal_3095 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1700
  signal new_AGEMA_signal_3096 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1701
  signal new_AGEMA_signal_3097 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1702
  signal new_AGEMA_signal_3098 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1703
  signal new_AGEMA_signal_3099 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1704
  signal new_AGEMA_signal_3100 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1705
  signal new_AGEMA_signal_3101 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1706
  signal new_AGEMA_signal_3102 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1707
  signal new_AGEMA_signal_3103 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1708
  signal new_AGEMA_signal_3104 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1709
  signal new_AGEMA_signal_3105 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1710
  signal new_AGEMA_signal_3106 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1711
  signal new_AGEMA_signal_3107 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1712
  signal new_AGEMA_signal_3108 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1713
  signal new_AGEMA_signal_3109 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1714
  signal new_AGEMA_signal_3110 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1715
  signal new_AGEMA_signal_3111 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1716
  signal new_AGEMA_signal_3112 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1717
  signal new_AGEMA_signal_3113 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1718
  signal new_AGEMA_signal_3114 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1719
  signal new_AGEMA_signal_3115 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1720
  signal new_AGEMA_signal_3116 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1721
  signal new_AGEMA_signal_3117 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1722
  signal new_AGEMA_signal_3118 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1723
  signal new_AGEMA_signal_3119 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1724
  signal new_AGEMA_signal_3120 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1725
  signal new_AGEMA_signal_3121 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1726
  signal new_AGEMA_signal_3122 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1727
  signal new_AGEMA_signal_3123 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1728
  signal new_AGEMA_signal_3124 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1729
  signal new_AGEMA_signal_3125 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1730
  signal new_AGEMA_signal_3126 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1731
  signal new_AGEMA_signal_3127 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1732
  signal new_AGEMA_signal_3128 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1733
  signal new_AGEMA_signal_3129 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1734
  signal new_AGEMA_signal_3130 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1735
  signal new_AGEMA_signal_3131 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1736
  signal new_AGEMA_signal_3132 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1737
  signal new_AGEMA_signal_3133 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1738
  signal new_AGEMA_signal_3134 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1739
  signal new_AGEMA_signal_3135 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1740
  signal new_AGEMA_signal_3136 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1741
  signal new_AGEMA_signal_3137 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1742
  signal new_AGEMA_signal_3138 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1743
  signal new_AGEMA_signal_3139 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1744
  signal new_AGEMA_signal_3140 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1745
  signal new_AGEMA_signal_3141 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1746
  signal new_AGEMA_signal_3142 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1747
  signal new_AGEMA_signal_3143 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1748
  signal new_AGEMA_signal_3144 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1749
  signal new_AGEMA_signal_3145 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1750
  signal new_AGEMA_signal_3146 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1751
  signal new_AGEMA_signal_3147 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1752
  signal new_AGEMA_signal_3148 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1753
  signal new_AGEMA_signal_3149 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1754
  signal new_AGEMA_signal_3150 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1755
  signal new_AGEMA_signal_3151 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1756
  signal new_AGEMA_signal_3152 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1757
  signal new_AGEMA_signal_3153 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1758
  signal new_AGEMA_signal_3154 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1759
  signal new_AGEMA_signal_3155 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1760
  signal new_AGEMA_signal_3156 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1761
  signal new_AGEMA_signal_3157 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1762
  signal new_AGEMA_signal_3158 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1763
  signal new_AGEMA_signal_3159 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1764
  signal new_AGEMA_signal_3160 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1765
  signal new_AGEMA_signal_3161 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1766
  signal new_AGEMA_signal_3162 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1767
  signal new_AGEMA_signal_3163 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1768
  signal new_AGEMA_signal_3164 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1769
  signal new_AGEMA_signal_3165 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1770
  signal new_AGEMA_signal_3166 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1771
  signal new_AGEMA_signal_3167 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1772
  signal new_AGEMA_signal_3168 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1773
  signal new_AGEMA_signal_3169 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1774
  signal new_AGEMA_signal_3170 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1775
  signal new_AGEMA_signal_3171 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1776
  signal new_AGEMA_signal_3172 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1777
  signal new_AGEMA_signal_3173 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1778
  signal new_AGEMA_signal_3174 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1779
  signal new_AGEMA_signal_3175 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1780
  signal new_AGEMA_signal_3176 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1781
  signal new_AGEMA_signal_3177 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1782
  signal new_AGEMA_signal_3178 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1783
  signal new_AGEMA_signal_3179 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1784
  signal new_AGEMA_signal_3180 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1785
  signal new_AGEMA_signal_3181 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1786
  signal new_AGEMA_signal_3182 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1787
  signal new_AGEMA_signal_3183 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1788
  signal new_AGEMA_signal_3184 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1789
  signal new_AGEMA_signal_3185 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1790
  signal new_AGEMA_signal_3186 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1791
  signal new_AGEMA_signal_3187 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1792
  signal new_AGEMA_signal_3188 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1793
  signal new_AGEMA_signal_3189 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1794
  signal new_AGEMA_signal_3190 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1795
  signal new_AGEMA_signal_3191 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1796
  signal new_AGEMA_signal_3192 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1797
  signal new_AGEMA_signal_3193 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1798
  signal new_AGEMA_signal_3194 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1799
  signal new_AGEMA_signal_3195 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1800
  signal new_AGEMA_signal_3196 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1801
  signal new_AGEMA_signal_3197 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1802
  signal new_AGEMA_signal_3198 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1803
  signal new_AGEMA_signal_3199 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1804
  signal new_AGEMA_signal_3200 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1805
  signal new_AGEMA_signal_3201 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1806
  signal new_AGEMA_signal_3202 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1807
  signal new_AGEMA_signal_3203 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1808
  signal new_AGEMA_signal_3204 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1809
  signal new_AGEMA_signal_3205 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1810
  signal new_AGEMA_signal_3206 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1811
  signal new_AGEMA_signal_3207 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1812
  signal new_AGEMA_signal_3208 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1813
  signal new_AGEMA_signal_3209 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1814
  signal new_AGEMA_signal_3210 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1815
  signal new_AGEMA_signal_3211 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1816
  signal new_AGEMA_signal_3212 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1817
  signal new_AGEMA_signal_3213 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1818
  signal new_AGEMA_signal_3214 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1819
  signal new_AGEMA_signal_3215 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1820
  signal new_AGEMA_signal_3216 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1821
  signal new_AGEMA_signal_3217 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1822
  signal new_AGEMA_signal_3218 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1823
  signal new_AGEMA_signal_3219 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1824
  signal new_AGEMA_signal_3220 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1825
  signal new_AGEMA_signal_3221 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1826
  signal new_AGEMA_signal_3222 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1827
  signal new_AGEMA_signal_3223 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1828
  signal new_AGEMA_signal_3224 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1829
  signal new_AGEMA_signal_3225 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1830
  signal new_AGEMA_signal_3226 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1831
  signal new_AGEMA_signal_3227 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1832
  signal new_AGEMA_signal_3228 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1833
  signal new_AGEMA_signal_3229 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1834
  signal new_AGEMA_signal_3230 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1835
  signal new_AGEMA_signal_3231 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1836
  signal new_AGEMA_signal_3232 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1837
  signal new_AGEMA_signal_3233 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1838
  signal new_AGEMA_signal_3234 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1839
  signal new_AGEMA_signal_3235 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1840
  signal new_AGEMA_signal_3236 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1841
  signal new_AGEMA_signal_3237 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1842
  signal new_AGEMA_signal_3238 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1843
  signal new_AGEMA_signal_3239 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1844
  signal new_AGEMA_signal_3240 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1845
  signal new_AGEMA_signal_3241 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1846
  signal new_AGEMA_signal_3242 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1847
  signal new_AGEMA_signal_3243 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1848
  signal new_AGEMA_signal_3244 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1849
  signal new_AGEMA_signal_3245 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1850
  signal new_AGEMA_signal_3246 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1851
  signal new_AGEMA_signal_3247 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1852
  signal new_AGEMA_signal_3248 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1853
  signal new_AGEMA_signal_3249 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1854
  signal new_AGEMA_signal_3250 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1855
  signal new_AGEMA_signal_3251 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1856
  signal new_AGEMA_signal_3252 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1857
  signal new_AGEMA_signal_3253 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1858
  signal new_AGEMA_signal_3254 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1859
  signal new_AGEMA_signal_3255 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1860
  signal new_AGEMA_signal_3256 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1861
  signal new_AGEMA_signal_3257 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1862
  signal new_AGEMA_signal_3258 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1863
  signal new_AGEMA_signal_3259 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1864
  signal new_AGEMA_signal_3260 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1865
  signal new_AGEMA_signal_3261 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1866
  signal new_AGEMA_signal_3262 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1867
  signal new_AGEMA_signal_3263 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1868
  signal new_AGEMA_signal_3264 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1869
  signal new_AGEMA_signal_3265 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1870
  signal new_AGEMA_signal_3266 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1871
  signal new_AGEMA_signal_3267 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1872
  signal new_AGEMA_signal_3268 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1873
  signal new_AGEMA_signal_3269 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1874
  signal new_AGEMA_signal_3270 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1875
  signal new_AGEMA_signal_3271 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1876
  signal new_AGEMA_signal_3272 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1877
  signal new_AGEMA_signal_3273 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1878
  signal new_AGEMA_signal_3274 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1879
  signal new_AGEMA_signal_3275 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1880
  signal new_AGEMA_signal_3276 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1881
  signal new_AGEMA_signal_3277 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1882
  signal new_AGEMA_signal_3278 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1883
  signal new_AGEMA_signal_3279 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1884
  signal new_AGEMA_signal_3280 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1885
  signal new_AGEMA_signal_3281 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1886
  signal new_AGEMA_signal_3282 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1887
  signal new_AGEMA_signal_3283 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1888
  signal new_AGEMA_signal_3284 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1889
  signal new_AGEMA_signal_3285 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1890
  signal new_AGEMA_signal_3286 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1891
  signal new_AGEMA_signal_3287 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1892
  signal new_AGEMA_signal_3288 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1893
  signal new_AGEMA_signal_3289 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1894
  signal new_AGEMA_signal_3290 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1895
  signal new_AGEMA_signal_3291 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1896
  signal new_AGEMA_signal_3292 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1897
  signal new_AGEMA_signal_3293 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1898
  signal new_AGEMA_signal_3294 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1899
  signal new_AGEMA_signal_3295 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1900
  signal new_AGEMA_signal_3296 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1901
  signal new_AGEMA_signal_3297 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1902
  signal new_AGEMA_signal_3298 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1903
  signal new_AGEMA_signal_3299 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1904
  signal new_AGEMA_signal_3300 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1905
  signal new_AGEMA_signal_3301 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1906
  signal new_AGEMA_signal_3302 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1907
  signal new_AGEMA_signal_3303 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1908
  signal new_AGEMA_signal_3304 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1909
  signal new_AGEMA_signal_3305 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1910
  signal new_AGEMA_signal_3306 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1911
  signal new_AGEMA_signal_3307 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1912
  signal new_AGEMA_signal_3308 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1913
  signal new_AGEMA_signal_3309 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1914
  signal new_AGEMA_signal_3310 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1915
  signal new_AGEMA_signal_3311 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1916
  signal new_AGEMA_signal_3312 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1917
  signal new_AGEMA_signal_3313 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1918
  signal new_AGEMA_signal_3314 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1919
  signal new_AGEMA_signal_3315 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1920
  signal new_AGEMA_signal_3316 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1921
  signal new_AGEMA_signal_3317 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1922
  signal new_AGEMA_signal_3318 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1923
  signal new_AGEMA_signal_3319 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1924
  signal new_AGEMA_signal_3320 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1925
  signal new_AGEMA_signal_3321 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1926
  signal new_AGEMA_signal_3322 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1927
  signal new_AGEMA_signal_3323 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1928
  signal new_AGEMA_signal_3324 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1929
  signal new_AGEMA_signal_3325 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1930
  signal new_AGEMA_signal_3326 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1931
  signal new_AGEMA_signal_3327 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1932
  signal new_AGEMA_signal_3328 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1933
  signal new_AGEMA_signal_3329 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1934
  signal new_AGEMA_signal_3330 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1935
  signal new_AGEMA_signal_3331 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1936
  signal new_AGEMA_signal_3332 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1937
  signal new_AGEMA_signal_3333 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1938
  signal new_AGEMA_signal_3334 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1939
  signal new_AGEMA_signal_3335 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1940
  signal new_AGEMA_signal_3336 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1941
  signal new_AGEMA_signal_3337 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1942
  signal new_AGEMA_signal_3338 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1943
  signal new_AGEMA_signal_3339 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1944
  signal new_AGEMA_signal_3340 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1945
  signal new_AGEMA_signal_3341 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1946
  signal new_AGEMA_signal_3342 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1947
  signal new_AGEMA_signal_3343 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1948
  signal new_AGEMA_signal_3344 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1949
  signal new_AGEMA_signal_3345 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1950
  signal new_AGEMA_signal_3346 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1951
  signal new_AGEMA_signal_3347 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1952
  signal new_AGEMA_signal_3348 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1953
  signal new_AGEMA_signal_3349 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1954
  signal new_AGEMA_signal_3350 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1955
  signal new_AGEMA_signal_3351 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1956
  signal new_AGEMA_signal_3352 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1957
  signal new_AGEMA_signal_3353 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1958
  signal new_AGEMA_signal_3354 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1959
  signal new_AGEMA_signal_3355 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1960
  signal new_AGEMA_signal_3356 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1961
  signal new_AGEMA_signal_3357 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1962
  signal new_AGEMA_signal_3358 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1963
  signal new_AGEMA_signal_3359 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1964
  signal new_AGEMA_signal_3360 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1965
  signal new_AGEMA_signal_3361 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1966
  signal new_AGEMA_signal_3362 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1967
  signal new_AGEMA_signal_3363 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1968
  signal new_AGEMA_signal_3364 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1969
  signal new_AGEMA_signal_3365 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1970
  signal new_AGEMA_signal_3366 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1971
  signal new_AGEMA_signal_3367 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1972
  signal new_AGEMA_signal_3368 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1973
  signal new_AGEMA_signal_3369 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1974
  signal new_AGEMA_signal_3370 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1975
  signal new_AGEMA_signal_3371 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1976
  signal new_AGEMA_signal_3372 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1977
  signal new_AGEMA_signal_3373 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1978
  signal new_AGEMA_signal_3374 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1979
  signal new_AGEMA_signal_3375 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1980
  signal new_AGEMA_signal_3376 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1981
  signal new_AGEMA_signal_3377 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1982
  signal new_AGEMA_signal_3378 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1983
  signal new_AGEMA_signal_3379 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1984
  signal new_AGEMA_signal_3380 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1985
  signal new_AGEMA_signal_3381 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1986
  signal new_AGEMA_signal_3382 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1987
  signal new_AGEMA_signal_3383 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1988
  signal new_AGEMA_signal_3384 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1989
  signal new_AGEMA_signal_3385 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1990
  signal new_AGEMA_signal_3386 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1991
  signal new_AGEMA_signal_3387 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1992
  signal new_AGEMA_signal_3388 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1993
  signal new_AGEMA_signal_3389 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1994
  signal new_AGEMA_signal_3390 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1995
  signal new_AGEMA_signal_3391 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1996
  signal new_AGEMA_signal_3392 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1997
  signal new_AGEMA_signal_3393 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1998
  signal new_AGEMA_signal_3394 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1999
  signal new_AGEMA_signal_3395 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2000
  signal new_AGEMA_signal_3396 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2001
  signal new_AGEMA_signal_3397 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2002
  signal new_AGEMA_signal_3398 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2003
  signal new_AGEMA_signal_3399 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2004
  signal new_AGEMA_signal_3400 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2005
  signal new_AGEMA_signal_3401 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2006
  signal new_AGEMA_signal_3402 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2007
  signal new_AGEMA_signal_3403 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2008
  signal new_AGEMA_signal_3404 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2009
  signal new_AGEMA_signal_3405 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2010
  signal new_AGEMA_signal_3406 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2011
  signal new_AGEMA_signal_3407 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2012
  signal new_AGEMA_signal_3408 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2013
  signal new_AGEMA_signal_3409 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2014
  signal new_AGEMA_signal_3410 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2015
  signal new_AGEMA_signal_3411 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2016
  signal new_AGEMA_signal_3412 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2017
  signal new_AGEMA_signal_3413 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2018
  signal new_AGEMA_signal_3414 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2019
  signal new_AGEMA_signal_3415 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2020
  signal new_AGEMA_signal_3416 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2021
  signal new_AGEMA_signal_3417 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2022
  signal new_AGEMA_signal_3418 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2023
  signal new_AGEMA_signal_3419 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2024
  signal new_AGEMA_signal_3420 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2025
  signal new_AGEMA_signal_3421 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2026
  signal new_AGEMA_signal_3422 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2027
  signal new_AGEMA_signal_3423 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2028
  signal new_AGEMA_signal_3424 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2029
  signal new_AGEMA_signal_3425 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2030
  signal new_AGEMA_signal_3426 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2031
  signal new_AGEMA_signal_3427 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2032
  signal new_AGEMA_signal_3428 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2033
  signal new_AGEMA_signal_3429 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2034
  signal new_AGEMA_signal_3430 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2035
  signal new_AGEMA_signal_3431 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2036
  signal new_AGEMA_signal_3432 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2037
  signal new_AGEMA_signal_3433 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2038
  signal new_AGEMA_signal_3434 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2039
  signal new_AGEMA_signal_3435 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2040
  signal new_AGEMA_signal_3436 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2041
  signal new_AGEMA_signal_3437 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2042
  signal new_AGEMA_signal_3438 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2043
  signal new_AGEMA_signal_3439 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2044
  signal new_AGEMA_signal_3440 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2045
  signal new_AGEMA_signal_3441 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2046
  signal new_AGEMA_signal_3442 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2047
  signal new_AGEMA_signal_3443 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2048
  signal new_AGEMA_signal_3444 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2049
  signal new_AGEMA_signal_3445 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2050
  signal new_AGEMA_signal_3446 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2051
  signal new_AGEMA_signal_3447 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2052
  signal new_AGEMA_signal_3448 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2053
  signal new_AGEMA_signal_3449 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2054
  signal new_AGEMA_signal_3450 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2055
  signal new_AGEMA_signal_3451 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2056
  signal new_AGEMA_signal_3452 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2057
  signal new_AGEMA_signal_3453 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2058
  signal new_AGEMA_signal_3454 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2059
  signal new_AGEMA_signal_3455 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2060
  signal new_AGEMA_signal_3456 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2061
  signal new_AGEMA_signal_3457 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2062
  signal new_AGEMA_signal_3458 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2063
  signal new_AGEMA_signal_3459 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2064
  signal new_AGEMA_signal_3460 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2065
  signal new_AGEMA_signal_3461 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2066
  signal new_AGEMA_signal_3462 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2067
  signal new_AGEMA_signal_3463 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2068
  signal new_AGEMA_signal_3464 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2069
  signal new_AGEMA_signal_3465 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2070
  signal new_AGEMA_signal_3466 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2071
  signal new_AGEMA_signal_3467 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2072
  signal new_AGEMA_signal_3468 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2073
  signal new_AGEMA_signal_3469 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2074
  signal new_AGEMA_signal_3470 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2075
  signal new_AGEMA_signal_3471 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2076
  signal new_AGEMA_signal_3472 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2077
  signal new_AGEMA_signal_3473 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2078
  signal new_AGEMA_signal_3474 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2079
  signal new_AGEMA_signal_3475 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2080
  signal new_AGEMA_signal_3476 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2081
  signal new_AGEMA_signal_3477 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2082
  signal new_AGEMA_signal_3478 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2083
  signal new_AGEMA_signal_3479 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2084
  signal new_AGEMA_signal_3480 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2085
  signal new_AGEMA_signal_3481 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2086
  signal new_AGEMA_signal_3482 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2087
  signal new_AGEMA_signal_3483 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2088
  signal new_AGEMA_signal_3484 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2089
  signal new_AGEMA_signal_3485 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2090
  signal new_AGEMA_signal_3486 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2091
  signal new_AGEMA_signal_3487 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2092
  signal new_AGEMA_signal_3488 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2093
  signal new_AGEMA_signal_3489 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2094
  signal new_AGEMA_signal_3490 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2095
  signal new_AGEMA_signal_3491 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2096
  signal new_AGEMA_signal_3492 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2097
  signal new_AGEMA_signal_3493 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2098
  signal new_AGEMA_signal_3494 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2099
  signal new_AGEMA_signal_3495 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2100
  signal new_AGEMA_signal_3496 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2101
  signal new_AGEMA_signal_3497 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2102
  signal new_AGEMA_signal_3498 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2103
  signal new_AGEMA_signal_3499 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2104
  signal new_AGEMA_signal_3500 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2105
  signal new_AGEMA_signal_3501 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2106
  signal new_AGEMA_signal_3502 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2107
  signal new_AGEMA_signal_3503 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2108
  signal new_AGEMA_signal_3504 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2109
  signal new_AGEMA_signal_3505 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2110
  signal new_AGEMA_signal_3506 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2111
  signal new_AGEMA_signal_3507 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2112
  signal new_AGEMA_signal_3508 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2113
  signal new_AGEMA_signal_3509 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2114
  signal new_AGEMA_signal_3510 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2115
  signal new_AGEMA_signal_3511 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2116
  signal new_AGEMA_signal_3512 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2117
  signal new_AGEMA_signal_3513 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2118
  signal new_AGEMA_signal_3514 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2119
  signal new_AGEMA_signal_3515 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2120
  signal new_AGEMA_signal_3516 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2121
  signal new_AGEMA_signal_3517 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2122
  signal new_AGEMA_signal_3518 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2123
  signal new_AGEMA_signal_3519 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2124
  signal new_AGEMA_signal_3520 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2125
  signal new_AGEMA_signal_3521 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2126
  signal new_AGEMA_signal_3522 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2127
  signal new_AGEMA_signal_3523 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2128
  signal new_AGEMA_signal_3524 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2129
  signal new_AGEMA_signal_3525 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2130
  signal new_AGEMA_signal_3526 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2131
  signal new_AGEMA_signal_3527 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2132
  signal new_AGEMA_signal_3528 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2133
  signal new_AGEMA_signal_3529 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2134
  signal new_AGEMA_signal_3530 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2135
  signal new_AGEMA_signal_3531 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2136
  signal new_AGEMA_signal_3532 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2137
  signal new_AGEMA_signal_3533 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2138
  signal new_AGEMA_signal_3534 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2139
  signal new_AGEMA_signal_3535 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2140
  signal new_AGEMA_signal_3536 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2141
  signal new_AGEMA_signal_3537 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2142
  signal new_AGEMA_signal_3538 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2143
  signal new_AGEMA_signal_3539 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2144
  signal new_AGEMA_signal_3540 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2145
  signal new_AGEMA_signal_3541 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2146
  signal new_AGEMA_signal_3542 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2147
  signal new_AGEMA_signal_3543 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2148
  signal new_AGEMA_signal_3544 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2149
  signal new_AGEMA_signal_3545 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2150
  signal new_AGEMA_signal_3546 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2151
  signal new_AGEMA_signal_3547 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2152
  signal new_AGEMA_signal_3548 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2153
  signal new_AGEMA_signal_3549 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2154
  signal new_AGEMA_signal_3550 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2155
  signal new_AGEMA_signal_3551 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2156
  signal new_AGEMA_signal_3552 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2157
  signal new_AGEMA_signal_3553 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2158
  signal new_AGEMA_signal_3554 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2159
  signal new_AGEMA_signal_3555 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2160
  signal new_AGEMA_signal_3556 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2161
  signal new_AGEMA_signal_3557 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2162
  signal new_AGEMA_signal_3558 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2163
  signal new_AGEMA_signal_3559 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2164
  signal new_AGEMA_signal_3560 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2165
  signal new_AGEMA_signal_3561 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2166
  signal new_AGEMA_signal_3562 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2167
  signal new_AGEMA_signal_3563 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2168
  signal new_AGEMA_signal_3564 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2169
  signal new_AGEMA_signal_3565 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2170
  signal new_AGEMA_signal_3566 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2171
  signal new_AGEMA_signal_3567 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2172
  signal new_AGEMA_signal_3568 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2173
  signal new_AGEMA_signal_3569 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2174
  signal new_AGEMA_signal_3570 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2175
  signal new_AGEMA_signal_3571 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2176
  signal new_AGEMA_signal_3572 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2177
  signal new_AGEMA_signal_3573 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2178
  signal new_AGEMA_signal_3574 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2179
  signal new_AGEMA_signal_3575 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2180
  signal new_AGEMA_signal_3576 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2181
  signal new_AGEMA_signal_3577 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2182
  signal new_AGEMA_signal_3578 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2183
  signal new_AGEMA_signal_3579 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2184
  signal new_AGEMA_signal_3580 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2185
  signal new_AGEMA_signal_3581 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2186
  signal new_AGEMA_signal_3582 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2187
  signal new_AGEMA_signal_3583 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2188
  signal new_AGEMA_signal_3584 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2189
  signal new_AGEMA_signal_3585 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2190
  signal new_AGEMA_signal_3586 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2191
  signal new_AGEMA_signal_3587 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2192
  signal new_AGEMA_signal_3588 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2193
  signal new_AGEMA_signal_3589 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2194
  signal new_AGEMA_signal_3590 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2195
  signal new_AGEMA_signal_3591 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2196
  signal new_AGEMA_signal_3592 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2197
  signal new_AGEMA_signal_3593 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2198
  signal new_AGEMA_signal_3594 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2199
  signal new_AGEMA_signal_3595 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2200
  signal new_AGEMA_signal_3596 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2201
  signal new_AGEMA_signal_3597 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2202
  signal new_AGEMA_signal_3598 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2203
  signal new_AGEMA_signal_3599 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2204
  signal new_AGEMA_signal_3600 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2205
  signal new_AGEMA_signal_3601 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2206
  signal new_AGEMA_signal_3602 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2207
  signal new_AGEMA_signal_3603 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2208
  signal new_AGEMA_signal_3604 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2209
  signal new_AGEMA_signal_3605 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2210
  signal new_AGEMA_signal_3606 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2211
  signal new_AGEMA_signal_3607 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2212
  signal new_AGEMA_signal_3608 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2213
  signal new_AGEMA_signal_3609 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2214
  signal new_AGEMA_signal_3610 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2215
  signal new_AGEMA_signal_3611 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2216
  signal new_AGEMA_signal_3612 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2217
  signal new_AGEMA_signal_3613 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2218
  signal new_AGEMA_signal_3614 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2219
  signal new_AGEMA_signal_3615 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2220
  signal new_AGEMA_signal_3616 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2221
  signal new_AGEMA_signal_3617 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2222
  signal new_AGEMA_signal_3618 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2223
  signal new_AGEMA_signal_3619 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2224
  signal new_AGEMA_signal_3620 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2225
  signal new_AGEMA_signal_3621 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2226
  signal new_AGEMA_signal_3622 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2227
  signal new_AGEMA_signal_3623 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2228
  signal new_AGEMA_signal_3624 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2229
  signal new_AGEMA_signal_3625 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2230
  signal new_AGEMA_signal_3626 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2231
  signal new_AGEMA_signal_3627 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2232
  signal new_AGEMA_signal_3628 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2233
  signal new_AGEMA_signal_3629 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2234
  signal new_AGEMA_signal_3630 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2235
  signal new_AGEMA_signal_3631 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2236
  signal new_AGEMA_signal_3632 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2237
  signal new_AGEMA_signal_3633 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2238
  signal new_AGEMA_signal_3634 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2239
  signal new_AGEMA_signal_3635 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2240
  signal new_AGEMA_signal_3636 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2241
  signal new_AGEMA_signal_3637 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2242
  signal new_AGEMA_signal_3638 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2243
  signal new_AGEMA_signal_3639 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2244
  signal new_AGEMA_signal_3640 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2245
  signal new_AGEMA_signal_3641 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2246
  signal new_AGEMA_signal_3642 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2247
  signal new_AGEMA_signal_3643 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2248
  signal new_AGEMA_signal_3644 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2249
  signal new_AGEMA_signal_3645 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2250
  signal new_AGEMA_signal_3646 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2251
  signal new_AGEMA_signal_3647 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2252
  signal new_AGEMA_signal_3648 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2253
  signal new_AGEMA_signal_3649 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2254
  signal new_AGEMA_signal_3650 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2255
  signal new_AGEMA_signal_3651 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2256
  signal new_AGEMA_signal_3652 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2257
  signal new_AGEMA_signal_3653 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2258
  signal new_AGEMA_signal_3654 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2259
  signal new_AGEMA_signal_3655 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2260
  signal new_AGEMA_signal_3656 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2261
  signal new_AGEMA_signal_3657 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2262
  signal new_AGEMA_signal_3658 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2263
  signal new_AGEMA_signal_3659 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2264
  signal new_AGEMA_signal_3660 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2265
  signal new_AGEMA_signal_3661 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2266
  signal new_AGEMA_signal_3662 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2267
  signal new_AGEMA_signal_3663 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2268
  signal new_AGEMA_signal_3664 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2269
  signal new_AGEMA_signal_3665 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2270
  signal new_AGEMA_signal_3666 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2271
  signal new_AGEMA_signal_3667 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2272
  signal new_AGEMA_signal_3668 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2273
  signal new_AGEMA_signal_3669 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2274
  signal new_AGEMA_signal_3670 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2275
  signal new_AGEMA_signal_3671 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2276
  signal new_AGEMA_signal_3672 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2277
  signal new_AGEMA_signal_3673 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2278
  signal new_AGEMA_signal_3674 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2279
  signal new_AGEMA_signal_3675 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2280
  signal new_AGEMA_signal_3676 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2281
  signal new_AGEMA_signal_3677 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2282
  signal new_AGEMA_signal_3678 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2283
  signal new_AGEMA_signal_3679 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2284
  signal new_AGEMA_signal_3680 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2285
  signal new_AGEMA_signal_3681 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2286
  signal new_AGEMA_signal_3682 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2287
  signal new_AGEMA_signal_3683 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2288
  signal new_AGEMA_signal_3684 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2289
  signal new_AGEMA_signal_3685 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2290
  signal new_AGEMA_signal_3686 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2291
  signal new_AGEMA_signal_3687 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2292
  signal new_AGEMA_signal_3688 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2293
  signal new_AGEMA_signal_3689 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2294
  signal new_AGEMA_signal_3690 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2295
  signal new_AGEMA_signal_3691 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2296
  signal new_AGEMA_signal_3692 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2297
  signal new_AGEMA_signal_3693 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2298
  signal new_AGEMA_signal_3694 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2299
  signal new_AGEMA_signal_3695 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2300
  signal new_AGEMA_signal_3696 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2301
  signal new_AGEMA_signal_3697 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2302
  signal new_AGEMA_signal_3698 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2303
  signal new_AGEMA_signal_3699 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2304
  signal new_AGEMA_signal_3700 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2305
  signal new_AGEMA_signal_3701 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2306
  signal new_AGEMA_signal_3702 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2307
  signal new_AGEMA_signal_3703 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2308
  signal new_AGEMA_signal_3704 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2309
  signal new_AGEMA_signal_3705 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2310
  signal new_AGEMA_signal_3706 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2311
  signal new_AGEMA_signal_3707 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2312
  signal new_AGEMA_signal_3708 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2313
  signal new_AGEMA_signal_3709 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2314
  signal new_AGEMA_signal_3710 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2315
  signal new_AGEMA_signal_3711 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2316
  signal new_AGEMA_signal_3712 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2317
  signal new_AGEMA_signal_3713 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2318
  signal new_AGEMA_signal_3714 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2319
  signal new_AGEMA_signal_3715 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2320
  signal new_AGEMA_signal_3716 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2321
  signal new_AGEMA_signal_3717 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2322
  signal new_AGEMA_signal_3718 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2323
  signal new_AGEMA_signal_3719 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2324
  signal new_AGEMA_signal_3720 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2325
  signal new_AGEMA_signal_3721 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2326
  signal new_AGEMA_signal_3722 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2327
  signal new_AGEMA_signal_3723 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2328
  signal new_AGEMA_signal_3724 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2329
  signal new_AGEMA_signal_3725 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2330
  signal new_AGEMA_signal_3726 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2331
  signal new_AGEMA_signal_3727 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2332
  signal new_AGEMA_signal_3728 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2333
  signal new_AGEMA_signal_3729 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2334
  signal new_AGEMA_signal_3730 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2335
  signal new_AGEMA_signal_3731 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2336
  signal new_AGEMA_signal_3732 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2337
  signal new_AGEMA_signal_3733 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2338
  signal new_AGEMA_signal_3734 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2339
  signal new_AGEMA_signal_3735 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2340
  signal new_AGEMA_signal_3736 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2341
  signal new_AGEMA_signal_3737 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2342
  signal new_AGEMA_signal_3738 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2343
  signal new_AGEMA_signal_3739 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2344
  signal new_AGEMA_signal_3740 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2345
  signal new_AGEMA_signal_3741 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2346
  signal new_AGEMA_signal_3742 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2347
  signal new_AGEMA_signal_3743 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2348
  signal new_AGEMA_signal_3744 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2349
  signal new_AGEMA_signal_3745 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2350
  signal new_AGEMA_signal_3746 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2351
  signal new_AGEMA_signal_3747 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2352
  signal new_AGEMA_signal_3748 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2353
  signal new_AGEMA_signal_3749 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2354
  signal new_AGEMA_signal_3750 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2355
  signal new_AGEMA_signal_3751 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2356
  signal new_AGEMA_signal_3752 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2357
  signal new_AGEMA_signal_3753 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2358
  signal new_AGEMA_signal_3754 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2359
  signal new_AGEMA_signal_3755 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2360
  signal new_AGEMA_signal_3756 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2361
  signal new_AGEMA_signal_3757 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2362
  signal new_AGEMA_signal_3758 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2363
  signal new_AGEMA_signal_3759 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2364
  signal new_AGEMA_signal_3760 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2365
  signal new_AGEMA_signal_3761 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2366
  signal new_AGEMA_signal_3762 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2367
  signal new_AGEMA_signal_3763 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2368
  signal new_AGEMA_signal_3764 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2369
  signal new_AGEMA_signal_3765 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2370
  signal new_AGEMA_signal_3766 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2371
  signal new_AGEMA_signal_3767 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2372
  signal new_AGEMA_signal_3768 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2373
  signal new_AGEMA_signal_3769 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2374
  signal new_AGEMA_signal_3770 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2375
  signal new_AGEMA_signal_3771 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2376
  signal new_AGEMA_signal_3772 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2377
  signal new_AGEMA_signal_3773 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2378
  signal new_AGEMA_signal_3774 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2379
  signal new_AGEMA_signal_3775 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2380
  signal new_AGEMA_signal_3776 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2381
  signal new_AGEMA_signal_3777 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2382
  signal new_AGEMA_signal_3778 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2383
  signal new_AGEMA_signal_3779 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2384
  signal new_AGEMA_signal_3780 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2385
  signal new_AGEMA_signal_3781 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2386
  signal new_AGEMA_signal_3782 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2387
  signal new_AGEMA_signal_3783 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2388
  signal new_AGEMA_signal_3784 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2389
  signal new_AGEMA_signal_3785 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2390
  signal new_AGEMA_signal_3786 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2391
  signal new_AGEMA_signal_3787 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2392
  signal new_AGEMA_signal_3788 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2393
  signal new_AGEMA_signal_3789 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2394
  signal new_AGEMA_signal_3790 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2395
  signal new_AGEMA_signal_3791 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2396
  signal new_AGEMA_signal_3792 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2397
  signal new_AGEMA_signal_3793 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2398
  signal new_AGEMA_signal_3794 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2399
  signal new_AGEMA_signal_3795 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2400
  signal new_AGEMA_signal_3796 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2401
  signal new_AGEMA_signal_3797 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2402
  signal new_AGEMA_signal_3798 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2403
  signal new_AGEMA_signal_3799 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2404
  signal new_AGEMA_signal_3800 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2405
  signal new_AGEMA_signal_3801 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2406
  signal new_AGEMA_signal_3802 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2407
  signal new_AGEMA_signal_3803 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2408
  signal new_AGEMA_signal_3804 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2409
  signal new_AGEMA_signal_3805 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2410
  signal new_AGEMA_signal_3806 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2411
  signal new_AGEMA_signal_3807 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2412
  signal new_AGEMA_signal_3808 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2413
  signal new_AGEMA_signal_3809 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2414
  signal new_AGEMA_signal_3810 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2415
  signal new_AGEMA_signal_3811 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2416
  signal new_AGEMA_signal_3812 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2417
  signal new_AGEMA_signal_3813 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2418
  signal new_AGEMA_signal_3814 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2419
  signal new_AGEMA_signal_3815 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2420
  signal new_AGEMA_signal_3816 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2421
  signal new_AGEMA_signal_3817 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2422
  signal new_AGEMA_signal_3818 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2423
  signal new_AGEMA_signal_3819 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2424
  signal new_AGEMA_signal_3820 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2425
  signal new_AGEMA_signal_3821 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2426
  signal new_AGEMA_signal_3822 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2427
  signal new_AGEMA_signal_3823 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2428
  signal new_AGEMA_signal_3824 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2429
  signal new_AGEMA_signal_3825 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2430
  signal new_AGEMA_signal_3826 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2431
  signal new_AGEMA_signal_3827 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2432
  signal new_AGEMA_signal_3828 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2433
  signal new_AGEMA_signal_3829 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2434
  signal new_AGEMA_signal_3830 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2435
  signal new_AGEMA_signal_3831 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2436
  signal new_AGEMA_signal_3832 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2437
  signal new_AGEMA_signal_3833 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2438
  signal new_AGEMA_signal_3834 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2439
  signal new_AGEMA_signal_3835 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2440
  signal new_AGEMA_signal_3836 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2441
  signal new_AGEMA_signal_3837 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2442
  signal new_AGEMA_signal_3838 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2443
  signal new_AGEMA_signal_3839 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2444
  signal new_AGEMA_signal_3840 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2445
  signal new_AGEMA_signal_3841 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2446
  signal new_AGEMA_signal_3842 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2447
  signal new_AGEMA_signal_3843 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2448
  signal new_AGEMA_signal_3844 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2449
  signal new_AGEMA_signal_3845 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2450
  signal new_AGEMA_signal_3846 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2451
  signal new_AGEMA_signal_3847 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2452
  signal new_AGEMA_signal_3848 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2453
  signal new_AGEMA_signal_3849 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2454
  signal new_AGEMA_signal_3850 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2455
  signal new_AGEMA_signal_3851 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2456
  signal new_AGEMA_signal_3852 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2457
  signal new_AGEMA_signal_3853 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2458
  signal new_AGEMA_signal_3854 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2459
  signal new_AGEMA_signal_3855 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2460
  signal new_AGEMA_signal_3856 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2461
  signal new_AGEMA_signal_3857 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2462
  signal new_AGEMA_signal_3858 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2463
  signal new_AGEMA_signal_3859 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2464
  signal new_AGEMA_signal_3860 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2465
  signal new_AGEMA_signal_3861 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2466
  signal new_AGEMA_signal_3862 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2467
  signal new_AGEMA_signal_3863 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2468
  signal new_AGEMA_signal_3864 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2469
  signal new_AGEMA_signal_3865 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2470
  signal new_AGEMA_signal_3866 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2471
  signal new_AGEMA_signal_3867 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2472
  signal new_AGEMA_signal_3868 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2473
  signal new_AGEMA_signal_3869 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2474
  signal new_AGEMA_signal_3870 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2475
  signal new_AGEMA_signal_3871 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2476
  signal new_AGEMA_signal_3872 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2477
  signal new_AGEMA_signal_3873 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2478
  signal new_AGEMA_signal_3874 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2479
  signal new_AGEMA_signal_3875 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2480
  signal new_AGEMA_signal_3876 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2481
  signal new_AGEMA_signal_3877 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2482
  signal new_AGEMA_signal_3878 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2483
  signal new_AGEMA_signal_3879 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2484
  signal new_AGEMA_signal_3880 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2485
  signal new_AGEMA_signal_3881 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2486
  signal new_AGEMA_signal_3882 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2487
  signal new_AGEMA_signal_3883 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2488
  signal new_AGEMA_signal_3884 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2489
  signal new_AGEMA_signal_3885 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2490
  signal new_AGEMA_signal_3886 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2491
  signal new_AGEMA_signal_3887 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2492
  signal new_AGEMA_signal_3888 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2493
  signal new_AGEMA_signal_3889 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2494
  signal new_AGEMA_signal_3890 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2495
  signal new_AGEMA_signal_3891 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2496
  signal new_AGEMA_signal_3892 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2497
  signal new_AGEMA_signal_3893 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2498
  signal new_AGEMA_signal_3894 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2499
  signal new_AGEMA_signal_3895 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2500
  signal new_AGEMA_signal_3896 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2501
  signal new_AGEMA_signal_3897 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2502
  signal new_AGEMA_signal_3898 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2503
  signal new_AGEMA_signal_3899 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2504
  signal new_AGEMA_signal_3900 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2505
  signal new_AGEMA_signal_3901 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2506
  signal new_AGEMA_signal_3902 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2507
  signal new_AGEMA_signal_3903 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2508
  signal new_AGEMA_signal_3904 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2509
  signal new_AGEMA_signal_3905 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2510
  signal new_AGEMA_signal_3906 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2511
  signal new_AGEMA_signal_3907 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2512
  signal new_AGEMA_signal_3908 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2513
  signal new_AGEMA_signal_3909 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2514
  signal new_AGEMA_signal_3910 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2515
  signal new_AGEMA_signal_3911 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2516
  signal new_AGEMA_signal_3912 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2517
  signal new_AGEMA_signal_3913 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2518
  signal new_AGEMA_signal_3914 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2519
  signal new_AGEMA_signal_3915 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2520
  signal new_AGEMA_signal_3916 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2521
  signal new_AGEMA_signal_3917 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2522
  signal new_AGEMA_signal_3918 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2523
  signal new_AGEMA_signal_3919 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2524
  signal new_AGEMA_signal_3920 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2525
  signal new_AGEMA_signal_3921 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2526
  signal new_AGEMA_signal_3922 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2527
  signal new_AGEMA_signal_3923 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2528
  signal new_AGEMA_signal_3924 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2529
  signal new_AGEMA_signal_3925 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2530
  signal new_AGEMA_signal_3926 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2531
  signal new_AGEMA_signal_3927 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2532
  signal new_AGEMA_signal_3928 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2533
  signal new_AGEMA_signal_3929 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2534
  signal new_AGEMA_signal_3930 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2535
  signal new_AGEMA_signal_3931 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2536
  signal new_AGEMA_signal_3932 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2537
  signal new_AGEMA_signal_3933 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2538
  signal new_AGEMA_signal_3934 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2539
  signal new_AGEMA_signal_3935 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2540
  signal new_AGEMA_signal_3936 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2541
  signal new_AGEMA_signal_3937 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2542
  signal new_AGEMA_signal_3938 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2543
  signal new_AGEMA_signal_3939 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2544
  signal new_AGEMA_signal_3940 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2545
  signal new_AGEMA_signal_3941 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2546
  signal new_AGEMA_signal_3942 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2547
  signal new_AGEMA_signal_3943 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2548
  signal new_AGEMA_signal_3944 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2549
  signal new_AGEMA_signal_3945 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2550
  signal new_AGEMA_signal_3946 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2551
  signal new_AGEMA_signal_3947 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2552
  signal new_AGEMA_signal_3948 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2553
  signal new_AGEMA_signal_3949 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2554
  signal new_AGEMA_signal_3950 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2555
  signal new_AGEMA_signal_3951 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2556
  signal new_AGEMA_signal_3952 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2557
  signal new_AGEMA_signal_3953 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2558
  signal new_AGEMA_signal_3954 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2559
  signal new_AGEMA_signal_3955 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2560
  signal new_AGEMA_signal_3956 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2561
  signal new_AGEMA_signal_3957 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2562
  signal new_AGEMA_signal_3958 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2563
  signal new_AGEMA_signal_3959 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2564
  signal new_AGEMA_signal_3960 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2565
  signal new_AGEMA_signal_3961 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2566
  signal new_AGEMA_signal_3962 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2567
  signal new_AGEMA_signal_3963 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2568
  signal new_AGEMA_signal_3964 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2569
  signal new_AGEMA_signal_3965 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2570
  signal new_AGEMA_signal_3966 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2571
  signal new_AGEMA_signal_3967 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2572
  signal new_AGEMA_signal_3968 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2573
  signal new_AGEMA_signal_3969 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2574
  signal new_AGEMA_signal_3970 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2575
  signal new_AGEMA_signal_3971 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2576
  signal new_AGEMA_signal_3972 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2577
  signal new_AGEMA_signal_3973 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2578
  signal new_AGEMA_signal_3974 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2579
  signal new_AGEMA_signal_3975 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2580
  signal new_AGEMA_signal_3976 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2581
  signal new_AGEMA_signal_3977 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2582
  signal new_AGEMA_signal_3978 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2583
  signal new_AGEMA_signal_3979 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2584
  signal new_AGEMA_signal_3980 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2585
  signal new_AGEMA_signal_3981 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2586
  signal new_AGEMA_signal_3982 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2587
  signal new_AGEMA_signal_3983 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2588
  signal new_AGEMA_signal_3984 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2589
  signal new_AGEMA_signal_3985 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2590
  signal new_AGEMA_signal_3986 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2591
  signal new_AGEMA_signal_3987 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2592
  signal new_AGEMA_signal_3988 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2593
  signal new_AGEMA_signal_3989 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2594
  signal new_AGEMA_signal_3990 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2595
  signal new_AGEMA_signal_3991 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2596
  signal new_AGEMA_signal_3992 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2597
  signal new_AGEMA_signal_3993 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2598
  signal new_AGEMA_signal_3994 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2599
  signal new_AGEMA_signal_3995 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2600
  signal new_AGEMA_signal_3996 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2601
  signal new_AGEMA_signal_3997 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2602
  signal new_AGEMA_signal_3998 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2603
  signal new_AGEMA_signal_3999 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2604
  signal new_AGEMA_signal_4000 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2605
  signal new_AGEMA_signal_4001 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2606
  signal new_AGEMA_signal_4002 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2607
  signal new_AGEMA_signal_4003 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2608
  signal new_AGEMA_signal_4004 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2609
  signal new_AGEMA_signal_4005 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2610
  signal new_AGEMA_signal_4006 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2611
  signal new_AGEMA_signal_4007 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2612
  signal new_AGEMA_signal_4008 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2613
  signal new_AGEMA_signal_4009 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2614
  signal new_AGEMA_signal_4010 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2615
  signal new_AGEMA_signal_4011 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2616
  signal new_AGEMA_signal_4012 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2617
  signal new_AGEMA_signal_4013 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2618
  signal new_AGEMA_signal_4014 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2619
  signal new_AGEMA_signal_4015 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2620
  signal new_AGEMA_signal_4016 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2621
  signal new_AGEMA_signal_4017 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2622
  signal new_AGEMA_signal_4018 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2623
  signal new_AGEMA_signal_4019 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2624
  signal new_AGEMA_signal_4020 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2625
  signal new_AGEMA_signal_4021 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2626
  signal new_AGEMA_signal_4022 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2627
  signal new_AGEMA_signal_4023 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2628
  signal new_AGEMA_signal_4024 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2629
  signal new_AGEMA_signal_4025 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2630
  signal new_AGEMA_signal_4026 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2631
  signal new_AGEMA_signal_4027 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2632
  signal new_AGEMA_signal_4028 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2633
  signal new_AGEMA_signal_4029 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2634
  signal new_AGEMA_signal_4030 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2635
  signal new_AGEMA_signal_4031 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2636
  signal new_AGEMA_signal_4032 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2637
  signal new_AGEMA_signal_4033 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2638
  signal new_AGEMA_signal_4034 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2639
  signal new_AGEMA_signal_4035 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2640
  signal new_AGEMA_signal_4036 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2641
  signal new_AGEMA_signal_4037 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2642
  signal new_AGEMA_signal_4038 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2643
  signal new_AGEMA_signal_4039 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2644
  signal new_AGEMA_signal_4040 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2645
  signal new_AGEMA_signal_4041 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2646
  signal new_AGEMA_signal_4042 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2647
  signal new_AGEMA_signal_4043 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2648
  signal new_AGEMA_signal_4044 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2649
  signal new_AGEMA_signal_4045 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2650
  signal new_AGEMA_signal_4046 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2651
  signal new_AGEMA_signal_4047 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2652
  signal new_AGEMA_signal_4048 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2653
  signal new_AGEMA_signal_4049 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2654
  signal new_AGEMA_signal_4050 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2655
  signal new_AGEMA_signal_4051 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2656
  signal new_AGEMA_signal_4052 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2657
  signal new_AGEMA_signal_4053 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2658
  signal new_AGEMA_signal_4054 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2659
  signal new_AGEMA_signal_4055 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2660
  signal new_AGEMA_signal_4056 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2661
  signal new_AGEMA_signal_4057 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2662
  signal new_AGEMA_signal_4058 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2663
  signal new_AGEMA_signal_4059 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2664
  signal new_AGEMA_signal_4060 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2665
  signal new_AGEMA_signal_4061 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2666
  signal new_AGEMA_signal_4062 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2667
  signal new_AGEMA_signal_4063 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2668
  signal new_AGEMA_signal_4064 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2669
  signal new_AGEMA_signal_4065 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2670
  signal new_AGEMA_signal_4066 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2671
  signal new_AGEMA_signal_4067 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2672
  signal new_AGEMA_signal_4068 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2673
  signal new_AGEMA_signal_4069 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2674
  signal new_AGEMA_signal_4070 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2675
  signal new_AGEMA_signal_4071 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2676
  signal new_AGEMA_signal_4072 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2677
  signal new_AGEMA_signal_4073 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2678
  signal new_AGEMA_signal_4074 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2679
  signal new_AGEMA_signal_4075 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2680
  signal new_AGEMA_signal_4076 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2681
  signal new_AGEMA_signal_4077 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2682
  signal new_AGEMA_signal_4078 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2683
  signal new_AGEMA_signal_4079 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2684
  signal new_AGEMA_signal_4080 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2685
  signal new_AGEMA_signal_4081 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2686
  signal new_AGEMA_signal_4082 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2687
  signal new_AGEMA_signal_4083 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2688
  signal new_AGEMA_signal_4084 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2689
  signal new_AGEMA_signal_4085 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2690
  signal new_AGEMA_signal_4086 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2691
  signal new_AGEMA_signal_4087 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2692
  signal new_AGEMA_signal_4088 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2693
  signal new_AGEMA_signal_4089 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2694
  signal new_AGEMA_signal_4090 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2695
  signal new_AGEMA_signal_4091 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2696
  signal new_AGEMA_signal_4092 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2697
  signal new_AGEMA_signal_4093 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2698
  signal new_AGEMA_signal_4094 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2699
  signal new_AGEMA_signal_4095 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2700
  signal new_AGEMA_signal_4096 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2701
  signal new_AGEMA_signal_4097 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2702
  signal new_AGEMA_signal_4098 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2703
  signal new_AGEMA_signal_4099 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2704
  signal new_AGEMA_signal_4100 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2705
  signal new_AGEMA_signal_4101 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2706
  signal new_AGEMA_signal_4102 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2707
  signal new_AGEMA_signal_4103 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2708
  signal new_AGEMA_signal_4104 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2709
  signal new_AGEMA_signal_4105 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2710
  signal new_AGEMA_signal_4106 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2711
  signal new_AGEMA_signal_4107 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2712
  signal new_AGEMA_signal_4108 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2713
  signal new_AGEMA_signal_4109 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2714
  signal new_AGEMA_signal_4110 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2715
  signal new_AGEMA_signal_4111 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2716
  signal new_AGEMA_signal_4112 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2717
  signal new_AGEMA_signal_4113 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2718
  signal new_AGEMA_signal_4114 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2719
  signal new_AGEMA_signal_4115 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2720
  signal new_AGEMA_signal_4116 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2721
  signal new_AGEMA_signal_4117 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2722
  signal new_AGEMA_signal_4118 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2723
  signal new_AGEMA_signal_4119 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2724
  signal new_AGEMA_signal_4120 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2725
  signal new_AGEMA_signal_4121 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2726
  signal new_AGEMA_signal_4122 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2727
  signal new_AGEMA_signal_4123 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2728
  signal new_AGEMA_signal_4124 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2729
  signal new_AGEMA_signal_4125 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2730
  signal new_AGEMA_signal_4126 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2731
  signal new_AGEMA_signal_4127 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2732
  signal new_AGEMA_signal_4128 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2733
  signal new_AGEMA_signal_4129 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2734
  signal new_AGEMA_signal_4130 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2735
  signal new_AGEMA_signal_4131 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2736
  signal new_AGEMA_signal_4132 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2737
  signal new_AGEMA_signal_4133 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2738
  signal new_AGEMA_signal_4134 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2739
  signal new_AGEMA_signal_4136 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2740
  signal new_AGEMA_signal_4137 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2741
  signal new_AGEMA_signal_4138 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2742
  signal new_AGEMA_signal_4140 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2743
  signal new_AGEMA_signal_4142 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2744
  signal new_AGEMA_signal_4143 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2745
  signal new_AGEMA_signal_4195 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2746
  signal new_AGEMA_signal_4197 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2747
  signal new_AGEMA_signal_4198 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2748
  signal new_AGEMA_signal_4199 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2749
  signal new_AGEMA_signal_4200 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2750
  signal new_AGEMA_signal_4201 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2751
  signal new_AGEMA_signal_4202 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2752
  signal new_AGEMA_signal_4203 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2753
  signal new_AGEMA_signal_4220 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2754
  signal new_AGEMA_signal_4221 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2755
  signal new_AGEMA_signal_4225 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2756
  signal new_AGEMA_signal_4226 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2757
  signal new_AGEMA_signal_4227 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2758
  signal new_AGEMA_signal_4230 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2759
  signal new_AGEMA_signal_4236 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2760
  signal new_AGEMA_signal_4237 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2761
  signal new_AGEMA_signal_4241 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2762
  signal new_AGEMA_signal_4242 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2763
  signal new_AGEMA_signal_4246 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2764
  signal new_AGEMA_signal_4248 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2765
  signal new_AGEMA_signal_4249 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2766
  signal new_AGEMA_signal_4252 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2767
  signal new_AGEMA_signal_4253 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2768
  signal new_AGEMA_signal_4254 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2769
  signal new_AGEMA_signal_4256 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2770
  signal new_AGEMA_signal_4257 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2771
  signal new_AGEMA_signal_4261 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2772
  signal new_AGEMA_signal_4262 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2773
  signal new_AGEMA_signal_4263 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2774
  signal new_AGEMA_signal_4264 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2775
  signal new_AGEMA_signal_4269 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2776
  signal new_AGEMA_signal_4271 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2777
  signal new_AGEMA_signal_4272 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2778
  signal new_AGEMA_signal_4276 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2779
  signal new_AGEMA_signal_4277 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2780
  signal new_AGEMA_signal_4278 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2781
  signal new_AGEMA_signal_4280 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2782
  signal new_AGEMA_signal_4284 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2783
  signal new_AGEMA_signal_4285 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2784
  signal new_AGEMA_signal_4287 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2785
  signal new_AGEMA_signal_4292 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2786
  signal new_AGEMA_signal_4293 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2787
  signal new_AGEMA_signal_4295 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2788
  signal new_AGEMA_signal_4296 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2789
  signal new_AGEMA_signal_4300 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2790
  signal new_AGEMA_signal_4302 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2791
  signal new_AGEMA_signal_4309 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2792
  signal new_AGEMA_signal_4310 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2793
  signal new_AGEMA_signal_4311 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2794
  signal new_AGEMA_signal_4313 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2795
  signal new_AGEMA_signal_4319 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2796
  signal new_AGEMA_signal_4320 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2797
  signal new_AGEMA_signal_4321 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2798
  signal new_AGEMA_signal_4322 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2799
  signal new_AGEMA_signal_4329 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2800
  signal new_AGEMA_signal_4330 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2801
  signal new_AGEMA_signal_4331 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2802
  signal new_AGEMA_signal_4332 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2803
  signal new_AGEMA_signal_4333 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2804
  signal new_AGEMA_signal_4334 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2805
  signal new_AGEMA_signal_4340 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2806
  signal new_AGEMA_signal_4341 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2807
  signal new_AGEMA_signal_4342 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2808
  signal new_AGEMA_signal_4343 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2809
  signal new_AGEMA_signal_4344 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2810
  signal new_AGEMA_signal_4345 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2811
  signal new_AGEMA_signal_4346 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2812
  signal new_AGEMA_signal_4347 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2813
  signal new_AGEMA_signal_4352 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2814
  signal new_AGEMA_signal_4355 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2815
  signal new_AGEMA_signal_4356 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2816
  signal new_AGEMA_signal_4357 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2817
  signal new_AGEMA_signal_4364 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2818
  signal new_AGEMA_signal_4365 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2819
  signal new_AGEMA_signal_4371 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2820
  signal new_AGEMA_signal_4372 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2821
  signal new_AGEMA_signal_4376 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2822
  signal new_AGEMA_signal_4377 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2823
  signal new_AGEMA_signal_4383 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2824
  signal new_AGEMA_signal_4384 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2825
  signal new_AGEMA_signal_4385 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2826
  signal new_AGEMA_signal_4386 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2827
  signal new_AGEMA_signal_4387 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2828
  signal new_AGEMA_signal_4388 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2829
  signal new_AGEMA_signal_4389 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2830
  signal new_AGEMA_signal_4390 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2831
  signal new_AGEMA_signal_4391 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2832
  signal new_AGEMA_signal_4392 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2833
  signal new_AGEMA_signal_4393 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2834
  signal new_AGEMA_signal_4394 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2835
  signal new_AGEMA_signal_4395 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2836
  signal new_AGEMA_signal_4396 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2837
  signal new_AGEMA_signal_4397 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2838
  signal new_AGEMA_signal_4398 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2839
  signal new_AGEMA_signal_4399 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2840
  signal new_AGEMA_signal_4400 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2841
  signal new_AGEMA_signal_4401 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2842
  signal new_AGEMA_signal_4402 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2843
  signal new_AGEMA_signal_4403 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2844
  signal new_AGEMA_signal_4404 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2845
  signal new_AGEMA_signal_4405 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2846
  signal new_AGEMA_signal_4406 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2847
  signal new_AGEMA_signal_4407 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2848
  signal new_AGEMA_signal_4408 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2849
  signal new_AGEMA_signal_4409 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2850
  signal new_AGEMA_signal_4410 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2851
  signal new_AGEMA_signal_4411 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2852
  signal new_AGEMA_signal_4412 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2853
  signal new_AGEMA_signal_4413 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2854
  signal new_AGEMA_signal_4414 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2855
  signal new_AGEMA_signal_4415 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2856
  signal new_AGEMA_signal_4416 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2857
  signal new_AGEMA_signal_4417 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2858
  signal new_AGEMA_signal_4418 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2859
  signal new_AGEMA_signal_4419 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2860
  signal new_AGEMA_signal_4420 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2861
  signal new_AGEMA_signal_4421 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2862
  signal new_AGEMA_signal_4422 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2863
  signal new_AGEMA_signal_4423 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2864
  signal new_AGEMA_signal_4424 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2865
  signal new_AGEMA_signal_4425 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2866
  signal new_AGEMA_signal_4426 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2867
  signal new_AGEMA_signal_4427 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2868
  signal new_AGEMA_signal_4428 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2869
  signal new_AGEMA_signal_4429 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2870
  signal new_AGEMA_signal_4430 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2871
  signal new_AGEMA_signal_4431 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2872
  signal new_AGEMA_signal_4432 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2873
  signal new_AGEMA_signal_4433 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2874
  signal new_AGEMA_signal_4434 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2875
  signal new_AGEMA_signal_4435 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2876
  signal new_AGEMA_signal_4436 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2877
  signal new_AGEMA_signal_4439 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2878
  signal new_AGEMA_signal_4441 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2879
  signal new_AGEMA_signal_4442 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2880
  signal new_AGEMA_signal_4443 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2881
  signal new_AGEMA_signal_4444 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2882
  signal new_AGEMA_signal_4445 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2883
  signal new_AGEMA_signal_4446 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2884
  signal new_AGEMA_signal_4447 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2885
  signal new_AGEMA_signal_4448 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2886
  signal new_AGEMA_signal_4449 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2887
  signal new_AGEMA_signal_4450 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2888
  signal new_AGEMA_signal_4451 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2889
  signal new_AGEMA_signal_4452 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2890
  signal new_AGEMA_signal_4496 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2891
  signal new_AGEMA_signal_4499 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2892
  signal new_AGEMA_signal_4500 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2893
  signal new_AGEMA_signal_4504 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2894
  signal new_AGEMA_signal_4505 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2895
  signal new_AGEMA_signal_4506 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2896
  signal new_AGEMA_signal_4510 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2897
  signal new_AGEMA_signal_4511 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2898
  signal new_AGEMA_signal_4550 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2899
  signal new_AGEMA_signal_4551 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2900
  signal new_AGEMA_signal_4558 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2901
  signal new_AGEMA_signal_4564 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2902
  signal new_AGEMA_signal_4565 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2903
  signal new_AGEMA_signal_4566 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2904
  signal new_AGEMA_signal_4570 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2905
  signal new_AGEMA_signal_4577 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2906
  signal new_AGEMA_signal_4578 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2907
  signal new_AGEMA_signal_4579 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2908
  signal new_AGEMA_signal_4580 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2909
  signal new_AGEMA_signal_4586 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2910
  signal new_AGEMA_signal_4591 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2911
  signal new_AGEMA_signal_4592 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2912
  signal new_AGEMA_signal_4593 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2913
  signal new_AGEMA_signal_4594 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2914
  signal new_AGEMA_signal_4596 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2915
  signal new_AGEMA_signal_4597 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2916
  signal new_AGEMA_signal_4598 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2917
  signal new_AGEMA_signal_4602 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2918
  signal new_AGEMA_signal_4603 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2919
  signal new_AGEMA_signal_4604 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2920
  signal new_AGEMA_signal_4605 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2921
  signal new_AGEMA_signal_4607 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2922
  signal new_AGEMA_signal_4608 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2923
  signal new_AGEMA_signal_4611 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2924
  signal new_AGEMA_signal_4614 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2925
  signal new_AGEMA_signal_4617 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2926
  signal new_AGEMA_signal_4618 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2927
  signal new_AGEMA_signal_4619 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2928
  signal new_AGEMA_signal_4621 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2929
  signal new_AGEMA_signal_4622 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2930
  signal new_AGEMA_signal_4627 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2931
  signal new_AGEMA_signal_4628 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2932
  signal new_AGEMA_signal_4639 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2933
  signal new_AGEMA_signal_4642 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2934
  signal new_AGEMA_signal_4643 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2935
  signal new_AGEMA_signal_4651 : std_logic;  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2936
  signal y0 : std_logic_vector(63 downto 0);  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1251
  signal y2 : std_logic_vector(1 downto 0);  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1252
  signal y4 : std_logic_vector(63 downto 0);  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1253
  signal z0 : std_logic_vector(63 downto 0);  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1254
  signal z1 : std_logic_vector(63 downto 0);  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1255
  signal z2 : std_logic_vector(63 downto 0);  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1256
  signal z3 : std_logic_vector(63 downto 0);  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1257
  signal z4 : std_logic_vector(63 downto 0);  -- Declared at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:1258
  signal LPM_q_ivl_7 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_47 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_57 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_65 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_76 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_86 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_94 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_105 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_115 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_123 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_134 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_144 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_152 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_163 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_173 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_181 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_192 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_202 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_210 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_221 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_231 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_239 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_250 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_260 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_268 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_279 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_289 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_297 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_308 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_318 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_326 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_337 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_347 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_355 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_366 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_376 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_384 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_395 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_405 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_413 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_424 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_434 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_442 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_453 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_463 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_471 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_482 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_492 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_500 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_511 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_521 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_529 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_540 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_550 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_558 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_569 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_579 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_587 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_598 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_608 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_616 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_627 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_637 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_645 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_656 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_666 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_674 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_685 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_695 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_703 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_714 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_724 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_732 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_743 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_753 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_761 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_772 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_782 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_790 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_801 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_811 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_819 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_830 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_840 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_848 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_859 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_869 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_877 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_888 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_898 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_906 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_917 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_927 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_935 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_946 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_956 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_964 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_975 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_985 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_993 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1004 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1014 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1022 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1033 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1043 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1051 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1062 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1072 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1080 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1091 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1101 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1109 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1120 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1130 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1138 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1149 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1159 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1167 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1178 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1188 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1196 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1207 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1217 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1225 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1236 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1246 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1254 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1265 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1275 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1283 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1294 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1304 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1312 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1323 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1333 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1341 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1352 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1362 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1370 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1381 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1391 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1399 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1410 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1420 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1428 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1439 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1449 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1457 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1468 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1478 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1486 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1497 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1507 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1515 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1526 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1536 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1544 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1555 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1565 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1573 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1584 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1594 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1602 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1613 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1623 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1631 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1642 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1652 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1660 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1671 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1681 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1689 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1700 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1710 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1718 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1729 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1739 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1747 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1758 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1768 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1776 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1787 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1797 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1805 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1816 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1826 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1834 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1845 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1855 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1863 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1874 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1884 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1892 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1903 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1913 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1921 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1932 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1942 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1950 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1961 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_1971 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1979 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_1990 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2000 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2008 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2019 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2029 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2037 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2048 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2058 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2066 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2077 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2087 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2095 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2106 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2116 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2124 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2135 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2145 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2153 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2164 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2174 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2182 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2193 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2203 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2211 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2222 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2232 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2240 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2251 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2261 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2269 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2280 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2290 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2298 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2309 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2319 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2327 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2338 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2348 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2356 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2367 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2377 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2385 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2396 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2406 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2414 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2425 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2435 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2443 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2454 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2464 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2472 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2483 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2493 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2501 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2512 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2522 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2530 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2541 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2551 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2559 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2570 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2580 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2588 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2599 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2609 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2617 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2628 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2638 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2646 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2657 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2667 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2675 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2686 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2696 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2704 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2715 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2725 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2733 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2744 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2754 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2762 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2773 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2783 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2791 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2802 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2812 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2820 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2831 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2841 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2849 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2860 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2870 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2878 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2889 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2899 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2907 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2918 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2928 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2936 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2947 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2957 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2965 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2976 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_2986 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_2994 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3005 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3015 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3023 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3034 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3044 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3052 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3063 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3073 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3081 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3092 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3102 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3110 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3121 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3131 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3139 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3150 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3160 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3168 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3179 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3189 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3197 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3208 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3218 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3226 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3237 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3247 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3255 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3266 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3276 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3284 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3295 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3305 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3313 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3324 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3334 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3342 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3353 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3363 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3371 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3382 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3392 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3400 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3411 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3421 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3429 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3440 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3450 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3458 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3469 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3479 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3487 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3498 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3508 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3516 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3527 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3537 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3545 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3556 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3566 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3574 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3585 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3595 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3603 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3614 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3624 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3632 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3643 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3653 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3661 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3672 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3682 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3690 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3701 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3711 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3719 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3730 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3738 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3746 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3757 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3765 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3773 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3784 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3792 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3800 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3811 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3819 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3827 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3838 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3846 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3854 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3865 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3873 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3881 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3892 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3900 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3908 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3919 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3927 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3935 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3946 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3954 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3962 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3973 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_3981 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_3989 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4000 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4008 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4016 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4027 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4035 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4043 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4054 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4062 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4070 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4081 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4089 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4097 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4108 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4116 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4124 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4135 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4143 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4151 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4162 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4170 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4178 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4189 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4197 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4205 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4216 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4224 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4232 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4243 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4251 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4259 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4270 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4278 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4286 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4297 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4305 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4313 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4324 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4332 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4340 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4351 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4359 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4367 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4378 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4386 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4394 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4405 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4413 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4421 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4432 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4440 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4448 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4459 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4467 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4475 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4486 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4494 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4502 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4513 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4521 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4529 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4540 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4548 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4556 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4567 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4575 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4583 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4594 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4602 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4610 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4621 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4629 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4637 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4648 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4656 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4664 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4675 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4683 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4691 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4702 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4710 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4718 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4729 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4737 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4745 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4756 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4764 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4772 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4783 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4791 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4799 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4810 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4818 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4826 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4837 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4845 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4853 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4864 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4872 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4880 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4891 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4899 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4907 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4918 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4926 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4934 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4945 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4953 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4961 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4972 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_4980 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4988 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_4999 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5007 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5015 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5026 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5034 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5042 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5053 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5061 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5069 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5080 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5088 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5096 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5107 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5115 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5123 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5134 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5142 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5150 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5161 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5169 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5177 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5188 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5196 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5204 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5215 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5223 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5231 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5242 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5250 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5258 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5269 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5277 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5285 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5296 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5304 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5312 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5323 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5331 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5339 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5350 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5358 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5366 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5377 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5385 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5393 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5404 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5412 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5420 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5431 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5439 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5447 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5458 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5466 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5474 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5485 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5493 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5501 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5512 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5520 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5528 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5539 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5547 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5555 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5566 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5574 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5582 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5593 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5601 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5602 : std_logic;
  signal LPM_q_ivl_5607 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5616 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5626 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5634 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5645 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5653 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5661 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5672 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5680 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5688 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5699 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5707 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5715 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5726 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5734 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5742 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5749 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5757 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5765 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5776 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5784 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5785 : std_logic;
  signal LPM_q_ivl_5787 : std_logic;
  signal LPM_q_ivl_5796 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5807 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5815 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5821 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5828 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5838 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5846 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5857 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5865 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5866 : std_logic;
  signal LPM_q_ivl_5871 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5880 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5888 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5889 : std_logic;
  signal LPM_q_ivl_5891 : std_logic;
  signal LPM_q_ivl_5898 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5909 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5917 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5925 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5932 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5940 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5946 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5957 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5965 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5969 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5980 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_5988 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_5996 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_6007 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_6015 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_6021 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_6028 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_6036 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_6044 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_6055 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_6063 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_6069 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_6076 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_6084 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_6088 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6090 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6095 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6097 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6102 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6104 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6109 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6111 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6116 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6118 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6123 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6125 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6130 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6132 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6137 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6139 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6144 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6146 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6151 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6153 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6158 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6160 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6165 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6167 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6172 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6174 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6179 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6181 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6186 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6188 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6193 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6195 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6200 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6202 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6207 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6209 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6214 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6216 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6221 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6223 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6228 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6230 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6235 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6237 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6242 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6244 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6249 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6251 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6256 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6258 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6263 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6265 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6270 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6272 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6277 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6279 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6284 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6286 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6291 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6293 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6298 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6300 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6305 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6307 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6312 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6314 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6319 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6321 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6326 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6328 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6333 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6335 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6340 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6342 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6347 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6349 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6354 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6356 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6361 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6363 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6368 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6370 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6375 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6377 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6382 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6384 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6389 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6391 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6396 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6398 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6403 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6405 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6410 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6412 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6417 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6419 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6424 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6426 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6431 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6433 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6438 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6440 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6445 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6447 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6452 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6454 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6459 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6461 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6466 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6468 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6473 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6475 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6480 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6482 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6487 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6489 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6494 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6496 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6501 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6503 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6508 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6510 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6515 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6517 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6522 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6524 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6529 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6531 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6538 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6540 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6547 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6549 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6556 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6558 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6565 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6567 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6574 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6576 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6583 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6585 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6592 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6594 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6601 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6603 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6610 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6612 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6619 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6621 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6628 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6630 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6637 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6639 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6646 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6648 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6655 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6657 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6664 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6666 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6673 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6675 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6682 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6684 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6691 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6693 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6700 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6702 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6709 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6711 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6718 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6720 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6727 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6729 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6736 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6738 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6745 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6747 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6754 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6756 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6763 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6765 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6772 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6774 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6781 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6783 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6790 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6792 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6799 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6801 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6808 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6810 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6817 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6819 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6826 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6828 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6835 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6837 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6844 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6846 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6853 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6855 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6862 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6864 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6871 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6873 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6880 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6882 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6889 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6891 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6898 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6900 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6907 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6909 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6916 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6918 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6925 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6927 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6934 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6936 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6943 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6945 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6952 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6954 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6961 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6963 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6970 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6972 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6979 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6981 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6988 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6990 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_6997 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_6999 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7006 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7008 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7015 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7017 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7024 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7026 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7033 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7035 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7042 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7044 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7051 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7053 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7060 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7062 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7069 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7071 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7078 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7080 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7087 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7089 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7096 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7098 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7105 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7107 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7114 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7116 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7123 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7125 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7132 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7134 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7141 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7143 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7150 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7152 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7159 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7161 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7168 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7170 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7177 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7179 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7186 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7188 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7195 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7197 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7204 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7206 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7213 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7215 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7222 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7224 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7231 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7233 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7240 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7242 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7249 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7251 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7258 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7260 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7267 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7269 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7276 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7278 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7285 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7287 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7294 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7296 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7303 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7305 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7312 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7314 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7321 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7323 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7330 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7332 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7339 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7341 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7348 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7350 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7357 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7359 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7366 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7368 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7375 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7377 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7384 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7386 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7393 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7395 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7402 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7404 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7411 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7413 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7420 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7422 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7429 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7431 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7438 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7440 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7447 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7449 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7456 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7458 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7465 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7467 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7474 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7476 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7483 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7485 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7492 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7494 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7501 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7503 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7510 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7512 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7519 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7521 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7528 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7530 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7537 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7539 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7546 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7548 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7555 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7557 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7564 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7566 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7573 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7575 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7582 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7584 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7591 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7593 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7600 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7602 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7609 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7611 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7618 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7620 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7627 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7629 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7636 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7638 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7645 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7647 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7654 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7656 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7663 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7665 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7672 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7674 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7681 : std_logic_vector(1 downto 0);
  signal LPM_d0_ivl_7683 : std_logic_vector(1 downto 0);
  signal LPM_q_ivl_7692 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7701 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7709 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7717 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7724 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7732 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7740 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7749 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7757 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7765 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7772 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7780 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7784 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7791 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7799 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7807 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7816 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7824 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7832 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7839 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7847 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7851 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7858 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7870 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7878 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7887 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7895 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7903 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7910 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7918 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7926 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7935 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7943 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7951 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7958 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7966 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7970 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7977 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_7985 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_7993 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8002 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8010 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8018 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8025 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8033 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8037 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8044 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8056 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8064 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8073 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8081 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8089 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8096 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8104 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8112 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8121 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8129 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8137 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8144 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8152 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8156 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8163 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8171 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8179 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8188 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8196 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8204 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8211 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8219 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8223 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8230 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8242 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8250 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8259 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8267 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8275 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8282 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8290 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8298 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8307 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8315 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8323 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8330 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8338 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8342 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8349 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8357 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8365 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8374 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8382 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8390 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8397 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8405 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8409 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8416 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8428 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8436 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8445 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8453 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8461 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8468 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8476 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8484 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8493 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8501 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8509 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8516 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8524 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8528 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8535 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8543 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8551 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8560 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8568 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8576 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8583 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8591 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8595 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8602 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8614 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8622 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8631 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8639 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8647 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8654 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8662 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8670 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8679 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8687 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8695 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8702 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8710 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8714 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8721 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8729 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8737 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8746 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8754 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8762 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8769 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8777 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8781 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8788 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8800 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8808 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8817 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8825 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8833 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8840 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8848 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8852 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8859 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8867 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8875 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8884 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8892 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8900 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8907 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8915 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8919 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8926 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8938 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8946 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8955 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8963 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8971 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8978 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_8986 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_8994 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9003 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9011 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9019 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9026 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9034 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9038 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9045 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9053 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9061 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9070 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9078 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9086 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9093 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9101 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9105 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9112 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9124 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9132 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9141 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9149 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9157 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9164 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9172 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9176 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9183 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9191 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9199 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9208 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9216 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9224 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9231 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9239 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9243 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9250 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9262 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9270 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9279 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9287 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9295 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9302 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9310 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9314 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9321 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9329 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9337 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9346 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9354 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9362 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9369 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9377 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9381 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9388 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9400 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9408 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9417 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9425 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9433 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9440 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9448 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9452 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9459 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9467 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9475 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9484 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9492 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9500 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9507 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9515 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9519 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9526 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9538 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9546 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9555 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9563 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9571 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9578 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9586 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9590 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9597 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9605 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9613 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9622 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9630 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9638 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9645 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9653 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9657 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9664 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9676 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9680 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9687 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9695 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9703 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9712 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9720 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9728 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9735 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9743 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9747 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9754 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9766 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9770 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9777 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9785 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9793 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9802 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9810 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9818 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9825 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9833 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9837 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9844 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9856 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9864 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9873 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9881 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9889 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9896 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9904 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9908 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9915 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9923 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9931 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9940 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9948 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9956 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9963 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9971 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9975 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_9982 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_9994 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10002 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10011 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10019 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10027 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10034 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10042 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10046 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10053 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10061 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10069 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10078 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10086 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10094 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10101 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10109 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10113 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10120 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10132 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10138 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10149 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10157 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10163 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10170 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10178 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10182 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10189 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10197 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10203 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10214 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10222 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10228 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10239 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10247 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10255 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10262 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10270 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10274 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10281 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10289 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10293 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10300 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10308 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10314 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10325 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10333 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10339 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10350 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10358 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10366 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10373 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10381 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10385 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10392 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10400 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10404 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10411 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10423 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10429 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10440 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10448 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10454 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10461 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10469 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10473 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10480 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10488 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10494 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10505 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10513 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10519 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10530 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10538 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10546 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10553 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10561 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10565 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10572 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10580 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10584 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10591 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10599 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10605 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10616 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10624 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10630 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10641 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10649 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10657 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10664 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10672 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10676 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10683 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10691 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10695 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10702 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10714 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10718 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10725 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10733 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10741 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10750 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10758 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10766 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10773 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10781 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10785 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10792 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10804 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10808 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10815 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10823 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10831 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10840 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10848 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10856 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10863 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10871 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10875 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10882 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10894 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10902 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10911 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10919 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10927 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10934 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10942 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10946 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10953 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10961 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10969 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10978 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_10986 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_10994 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11001 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11009 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11013 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11020 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11032 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11038 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11049 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11057 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11063 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11074 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11082 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11090 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11097 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11105 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11109 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11116 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11124 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11130 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11141 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11149 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11155 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11162 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11170 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11174 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11181 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11189 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11193 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11200 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11208 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11214 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11225 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11233 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11239 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11250 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11258 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11266 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11273 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11281 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11285 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11292 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11300 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11304 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11311 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11323 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11329 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11340 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11348 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11354 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11365 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11373 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11381 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11388 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11396 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11400 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11407 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11415 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11419 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11426 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11434 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11440 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11451 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11459 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11465 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11472 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11480 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11484 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11491 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11499 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11503 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11510 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11522 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11528 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11539 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11547 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11553 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11564 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11572 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11580 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11587 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11595 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11599 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11606 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11614 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11618 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11625 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11633 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11639 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11650 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11658 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11664 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11675 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11683 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11691 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11698 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11706 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11710 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11717 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11725 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11729 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11736 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11748 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11752 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11759 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11767 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11775 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11784 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11792 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11800 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11807 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11815 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11819 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11826 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11838 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11842 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11849 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11857 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11861 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11868 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11880 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11886 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11897 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11905 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11911 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11922 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11930 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11938 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11945 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11953 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11957 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11964 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11972 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11976 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11983 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_11991 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_11997 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12008 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12016 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12022 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12029 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12037 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12041 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12048 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12056 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12060 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12067 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12079 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12083 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12090 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12098 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12106 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12115 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12123 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12131 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12138 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12146 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12150 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12157 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12169 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12175 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12186 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12194 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12198 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12205 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12213 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12219 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12230 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12238 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12242 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12249 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12257 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12261 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12268 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12276 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12280 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12287 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12295 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12299 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12306 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12318 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12326 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12335 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12343 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12351 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12358 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12366 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12370 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12377 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12385 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12393 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12402 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12410 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12418 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12425 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12433 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12437 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12444 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12456 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12460 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12467 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12475 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12479 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12486 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12498 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12502 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12509 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12517 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12525 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12534 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12542 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12550 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12557 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12565 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12569 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12576 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12588 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12594 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12605 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12613 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12619 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12630 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12638 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12646 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12653 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12661 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12665 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12672 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12680 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12684 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12691 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12699 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12705 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12716 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12724 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12730 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12741 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12749 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12757 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12764 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12772 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12776 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12783 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12791 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12795 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12802 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12814 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12820 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12831 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12839 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12845 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12852 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12860 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12864 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12871 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12879 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12885 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12892 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12900 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12904 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12911 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12919 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12923 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12930 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12938 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12944 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12955 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12963 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12969 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12980 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_12988 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_12996 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13003 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13011 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13015 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13022 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13030 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13034 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13041 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13053 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13057 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13064 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13072 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13080 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13089 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13097 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13105 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13112 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13120 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13124 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13131 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13143 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13147 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13154 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13162 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13170 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13179 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13187 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13195 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13202 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13210 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13214 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13221 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13233 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13237 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13244 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13252 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13256 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13263 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13275 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13281 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13292 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13300 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13306 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13317 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13325 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13333 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13340 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13348 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13352 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13359 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13367 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13371 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13378 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13386 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13392 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13403 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13411 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13417 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13428 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13436 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13444 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13451 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13459 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13463 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13470 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13478 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13482 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13489 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13501 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13507 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13518 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13526 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13532 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13543 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13551 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13559 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13566 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13574 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13578 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13585 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13593 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13599 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13610 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13618 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13624 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13631 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13639 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13643 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13650 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13658 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13662 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13669 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13677 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13683 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13694 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13702 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13708 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13715 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13723 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13727 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13734 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13742 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13746 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13753 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13765 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13769 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13776 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13784 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13792 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13801 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13809 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13817 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13824 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13832 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13836 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13843 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13855 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13859 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13866 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13874 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13878 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13885 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13897 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13901 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13908 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13916 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13920 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13927 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13935 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13941 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13952 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13960 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13964 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13971 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_13979 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13983 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_13990 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14002 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14008 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14019 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14027 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14035 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14042 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14050 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14054 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14061 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14069 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14073 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14080 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14088 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14094 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14105 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14113 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14119 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14130 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14138 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14146 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14153 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14161 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14165 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14172 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14180 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14184 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14191 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14203 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14209 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14220 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14228 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14232 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14239 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14247 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14253 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14264 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14272 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14276 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14283 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14291 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14295 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14302 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14310 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14314 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14321 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14329 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14333 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14340 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14352 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14358 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14369 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14377 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14385 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14392 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14400 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14404 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14411 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14419 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14423 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14430 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14438 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14444 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14455 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14463 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14471 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14478 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14486 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14490 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14497 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14505 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14509 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14516 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14528 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14532 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14539 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14547 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14551 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14558 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14570 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14576 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14587 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14595 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14603 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14612 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14620 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14624 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14631 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14639 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14645 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14656 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14664 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14668 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14675 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14683 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14687 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14694 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14702 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14706 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14713 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14721 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14725 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14732 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14744 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14748 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14755 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14763 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14771 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14778 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14786 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14790 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14797 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14809 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14815 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14826 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14834 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14840 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14851 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14859 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14867 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14874 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14882 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14886 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14893 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14901 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14907 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14918 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14926 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14934 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14941 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14949 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14953 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14960 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14968 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14972 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14979 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_14987 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_14993 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15004 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15012 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15018 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15025 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15033 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15037 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15044 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15052 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15056 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15063 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15075 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15079 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15086 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15094 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15098 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15105 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15117 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15121 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15128 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15136 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15140 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15147 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15159 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15165 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15176 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15184 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15188 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15195 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15203 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15207 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15214 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15222 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15226 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15233 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15241 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15245 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15252 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15260 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15264 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15271 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15283 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15289 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15300 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15308 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15316 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15323 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15331 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15335 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15342 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15350 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15354 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15361 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15369 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15375 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15382 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15390 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15394 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15401 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15409 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15413 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15420 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15432 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15436 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15443 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15451 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15455 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15462 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15474 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15478 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15485 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15493 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15501 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15510 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15518 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15526 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15533 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15541 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15545 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15552 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15564 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15568 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15575 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15583 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15587 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15594 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15606 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15610 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15617 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15625 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15629 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15636 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15648 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15652 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15659 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15667 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15673 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15684 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15692 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15698 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15709 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15717 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15725 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15732 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15740 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15744 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15751 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15759 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15763 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15770 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15782 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15786 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15793 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15801 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15807 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15818 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15826 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15832 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15843 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15851 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15859 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15866 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15874 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15878 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15885 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15893 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15897 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15904 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15916 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15920 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15927 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15935 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15941 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15952 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15960 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15966 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15973 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_15981 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15985 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_15992 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16000 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16004 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16011 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16023 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16027 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16034 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16042 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16046 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16053 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16065 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16069 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16076 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16084 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16092 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16101 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16109 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16113 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16120 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16128 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16132 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16139 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16151 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16157 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16168 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16176 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16180 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16187 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16195 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16199 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16206 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16214 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16218 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16225 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16233 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16237 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16244 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16256 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16260 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16267 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16275 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16283 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16290 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16298 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16302 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16309 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16321 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16327 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16338 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16346 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16350 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16357 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16365 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16369 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16376 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16384 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16388 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16395 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16403 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16409 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16420 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16428 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16432 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16439 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16447 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16451 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16458 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16470 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16474 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16481 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16489 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16495 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16506 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16514 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16522 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16529 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16537 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16541 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16548 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16556 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16560 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16567 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16579 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16585 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16596 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16604 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16608 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16615 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16623 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16627 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16634 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16642 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16646 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16653 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16661 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16665 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16672 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16680 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16684 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16691 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16703 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16709 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16720 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16728 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16736 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16743 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16751 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16755 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16762 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16770 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16774 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16781 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16789 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16795 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16806 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16814 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16822 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16829 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16837 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16841 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16848 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16856 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16860 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16867 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16879 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16883 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16890 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16898 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16902 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16909 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16921 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16925 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16932 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16940 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16948 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16957 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16965 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16973 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16980 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_16988 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16992 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_16999 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17011 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17015 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17022 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17030 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17034 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17041 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17053 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17057 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17064 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17072 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17076 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17083 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17095 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17099 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17106 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17114 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17120 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17131 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17139 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17145 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17156 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17164 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17172 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17179 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17187 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17191 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17198 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17206 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17210 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17217 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17229 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17233 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17240 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17248 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17254 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17265 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17273 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17279 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17286 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17294 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17298 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17305 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17313 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17317 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17324 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17336 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17340 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17347 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17355 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17359 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17366 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17378 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17384 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17395 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17403 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17407 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17414 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17422 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17426 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17433 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17441 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17445 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17452 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17460 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17464 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17471 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17483 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17487 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17494 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17502 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17508 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17519 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17527 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17535 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17542 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17550 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17554 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17561 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17569 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17573 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17580 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17592 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17596 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17603 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17611 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17619 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17628 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17636 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17640 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17647 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17655 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17659 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17666 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17678 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17682 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17689 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17697 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17701 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17708 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17720 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17724 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17731 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17739 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17747 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17754 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17762 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17766 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17773 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17785 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17789 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17796 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17804 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17810 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17821 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17829 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17835 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17846 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17854 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17862 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17869 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17877 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17881 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17888 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17896 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17900 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17907 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17919 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17923 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17930 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17938 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17944 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17951 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17959 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17963 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17970 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_17978 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17982 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_17989 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18001 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18007 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18018 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18026 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18030 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18037 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18045 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18049 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18056 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18064 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18068 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18075 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18083 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18087 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18094 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18106 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18110 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18117 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18125 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18131 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18142 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18150 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18158 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18165 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18173 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18177 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18184 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18192 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18196 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18203 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18215 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18219 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18226 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18234 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18242 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18251 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18259 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18267 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18274 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18282 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18286 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18293 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18305 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18309 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18316 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18324 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18328 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18335 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18347 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18351 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18358 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18366 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18370 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18377 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18389 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18395 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18406 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18414 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18418 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18425 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18433 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18437 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18444 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18452 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18456 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18463 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18471 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18475 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18482 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18490 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18494 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18501 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18513 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18517 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18524 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18532 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18538 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18549 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18557 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18565 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18572 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18580 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18584 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18591 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18599 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18603 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18610 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18622 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18626 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18633 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18641 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18647 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18658 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18666 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18672 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18683 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18691 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18699 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18706 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18714 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18718 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18725 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18733 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18737 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18744 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18756 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18760 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18767 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18775 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18779 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18786 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18794 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18798 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18805 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18813 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18819 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18830 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18838 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18842 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18849 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18857 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18861 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18868 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18880 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18884 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18891 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18899 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18905 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18916 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18924 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18932 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18939 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18947 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18951 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18958 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18966 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18970 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18977 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_18989 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_18993 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19000 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19008 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19014 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19025 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19033 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19041 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19048 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19056 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19060 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19067 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19075 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19079 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19086 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19098 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19106 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19115 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19123 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19127 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19134 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19142 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19146 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19153 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19161 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19165 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19172 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19180 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19184 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19191 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19199 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19203 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19210 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19222 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19226 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19233 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19241 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19249 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19256 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19264 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19268 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19275 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19287 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19291 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19298 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19306 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19310 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19317 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19325 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19331 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19342 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19350 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19354 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19361 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19369 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19373 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19380 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19392 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19396 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19403 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19411 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19417 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19424 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19432 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19436 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19443 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19451 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19455 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19462 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19474 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19478 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19485 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19493 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19497 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19504 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19512 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19518 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19529 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19537 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19541 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19548 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19556 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19560 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19567 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19579 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19583 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19590 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19598 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19604 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19615 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19623 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19631 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19638 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19646 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19650 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19657 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19665 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19669 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19676 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19688 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19692 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19699 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19707 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19715 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19724 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19732 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19736 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19743 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19751 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19755 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19762 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19774 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19778 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19785 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19793 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19801 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19808 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19816 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19820 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19827 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19839 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19843 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19850 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19858 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19862 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19869 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19881 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19885 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19892 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19900 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19904 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19911 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19923 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19927 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19934 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19942 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19948 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19959 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19967 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19971 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19978 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_19986 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19990 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_19997 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20009 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20013 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20020 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20028 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20032 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20039 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20051 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20055 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20062 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20070 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20076 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20087 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20095 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20103 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20110 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20118 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20122 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20129 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20137 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20141 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20148 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20160 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20164 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20171 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20179 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20183 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20190 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20202 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20206 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20213 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20221 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20227 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20238 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20246 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20250 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20257 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20265 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20269 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20276 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20288 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20292 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20299 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20307 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20313 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20324 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20332 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20340 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20347 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20355 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20359 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20366 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20374 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20378 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20385 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20397 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20401 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20408 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20416 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20424 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20433 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20441 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20445 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20452 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20460 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20464 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20471 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20483 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20487 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20494 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20502 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20506 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20513 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20525 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20529 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20536 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20544 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20552 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20559 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20567 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20571 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20578 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20590 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20594 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20601 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20609 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20613 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20620 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20632 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20636 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20643 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20651 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20655 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20662 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20674 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20678 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20685 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20693 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20699 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20710 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20718 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20722 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20729 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20737 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20741 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20748 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20760 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20764 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20771 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20779 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20783 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20790 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20802 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20806 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20813 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20821 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20827 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20838 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20846 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20854 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20861 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20869 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20873 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20880 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20888 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20892 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20899 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20911 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20915 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20922 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20930 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20934 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20941 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20953 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20957 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20964 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20972 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20980 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_20989 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_20997 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21001 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21008 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21016 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21020 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21027 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21035 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21039 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21046 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21054 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21058 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21065 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21077 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21081 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21088 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21096 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21104 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21111 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21119 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21123 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21130 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21142 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21146 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21153 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21161 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21165 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21172 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21184 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21188 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21195 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21203 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21209 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21220 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21228 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21232 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21239 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21247 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21251 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21258 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21270 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21274 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21281 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21289 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21293 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21300 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21312 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21316 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21323 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21331 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21335 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21342 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21354 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21358 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21365 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21373 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21379 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21386 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21394 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21398 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21405 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21413 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21417 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21424 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21436 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21440 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21447 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21455 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21459 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21466 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21478 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21482 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21489 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21497 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21503 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21514 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21522 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21526 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21533 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21541 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21545 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21552 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21564 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21568 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21575 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21583 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21587 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21594 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21606 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21610 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21617 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21625 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21629 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21636 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21648 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21652 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21659 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21667 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21673 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21684 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21692 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21700 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21707 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21715 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21719 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21726 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21734 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21738 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21745 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21757 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21761 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21768 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21776 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21780 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21787 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21799 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21803 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21810 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21818 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21826 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21835 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21843 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21847 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21854 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21862 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21866 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21873 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21885 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21889 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21896 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21904 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21908 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21915 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21927 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21931 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21938 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21946 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21954 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21961 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21969 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21973 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21980 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_21992 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_21996 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22003 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22011 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22015 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22022 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22034 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22038 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22045 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22053 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22057 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22064 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22076 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22080 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22087 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22095 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22101 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22112 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22120 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22124 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22131 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22139 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22143 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22150 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22162 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22166 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22173 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22181 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22185 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22192 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22204 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22208 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22215 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22223 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22227 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22234 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22246 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22250 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22257 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22265 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22271 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22282 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22290 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22298 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22305 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22313 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22317 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22324 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22332 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22336 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22343 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22355 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22359 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22366 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22374 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22378 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22385 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22397 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22401 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22408 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22416 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22420 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22427 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22439 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22443 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22450 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22458 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22464 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22475 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22483 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22487 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22494 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22502 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22506 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22513 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22525 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22529 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22536 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22544 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22548 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22555 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22567 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22571 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22578 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22586 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22592 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22603 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22611 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22619 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22626 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22634 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22638 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22645 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22653 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22657 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22664 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22676 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22680 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22687 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22695 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22699 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22706 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22718 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22722 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22729 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22737 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22741 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22748 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22756 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22764 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22773 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22781 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22785 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22792 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22800 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22804 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22811 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22823 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22827 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22834 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22842 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22846 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22853 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22865 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22869 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22876 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22884 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22892 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22899 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22907 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22911 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22918 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22930 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22934 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22941 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22949 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22953 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22960 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22972 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22976 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22983 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_22991 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_22997 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23008 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23016 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23020 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23027 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23035 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23039 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23046 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23058 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23062 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23069 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23077 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23081 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23088 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23100 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23104 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23111 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23119 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23123 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23130 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23142 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23146 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23153 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23161 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23167 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23174 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23182 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23186 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23193 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23201 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23205 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23212 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23224 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23228 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23235 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23243 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23247 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23254 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23266 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23270 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23277 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23285 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23291 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23302 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23310 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23314 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23321 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23329 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23333 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23340 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23352 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23356 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23363 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23371 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23375 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23382 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23394 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23398 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23405 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23413 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23417 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23424 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23436 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23440 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23447 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23455 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23461 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23472 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23480 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23488 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23495 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23503 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23507 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23514 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23522 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23526 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23533 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23545 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23549 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23556 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23564 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23568 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23575 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23587 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23591 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23598 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23606 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23610 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23617 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23629 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23633 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23640 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23648 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23656 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23665 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23673 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23677 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23684 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23692 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23696 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23703 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23715 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23719 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23726 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23734 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23738 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23745 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23757 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23761 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23768 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23776 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23780 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23787 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23799 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23803 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23810 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23818 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23826 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23833 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23841 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23845 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23852 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23864 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23868 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23875 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23883 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23887 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23894 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23906 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23910 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23917 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23925 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23929 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23936 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23948 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23952 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23959 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23967 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23973 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23984 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_23992 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_23996 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24003 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24011 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24015 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24022 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24034 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24038 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24045 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24053 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24057 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24064 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24076 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24080 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24087 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24095 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24101 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24112 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24120 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24128 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24135 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24143 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24147 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24154 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24162 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24166 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24173 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24185 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24189 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24196 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24204 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24208 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24215 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24227 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24231 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24238 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24246 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24254 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24263 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24271 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24275 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24282 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24290 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24294 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24301 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24313 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24317 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24324 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24332 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24336 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24343 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24355 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24359 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24366 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24374 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24378 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24385 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24397 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24401 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24408 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24416 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24424 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24431 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24439 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24443 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24450 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24462 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24466 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24473 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24481 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24485 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24492 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24504 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24508 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24515 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24523 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24529 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24540 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24548 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24552 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24559 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24567 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24571 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24578 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24590 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24594 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24601 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24609 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24613 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24620 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24632 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24636 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24643 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24651 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24657 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24668 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24676 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24684 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24691 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24699 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24703 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24710 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24718 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24722 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24729 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24741 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24745 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24752 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24760 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24764 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24771 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24783 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24787 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24794 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24802 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24808 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24819 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24827 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24831 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24838 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24846 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24850 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24857 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24869 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24873 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24880 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24888 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24892 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24899 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24911 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24915 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24922 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24930 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24934 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24941 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24953 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24957 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24964 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24972 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24978 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_24989 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_24997 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25005 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25012 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25020 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25024 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25031 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25039 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25043 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25050 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25062 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25066 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25073 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25081 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25085 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25092 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25104 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25108 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25115 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25123 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25127 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25134 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25146 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25150 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25157 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25165 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25173 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25182 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25190 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25194 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25201 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25209 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25213 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25220 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25232 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25236 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25243 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25251 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25255 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25262 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25274 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25278 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25285 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25293 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25297 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25304 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25316 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25320 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25327 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25335 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25343 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25350 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25358 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25362 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25369 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25381 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25385 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25392 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25400 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25404 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25411 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25423 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25427 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25434 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25442 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25446 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25453 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25465 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25469 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25478 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25486 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25492 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25503 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25511 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25515 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25522 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25530 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25534 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25543 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25551 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25557 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25568 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25576 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25580 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25587 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25595 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25599 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25606 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25614 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25618 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25627 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25635 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25641 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25652 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25660 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25664 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25671 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25679 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25683 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25690 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25702 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25706 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25715 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25723 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25729 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25740 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25748 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25752 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25759 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25767 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25771 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25780 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25788 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25794 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25805 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25813 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25817 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25824 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25832 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25836 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25843 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25851 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25855 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25864 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25872 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25878 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25889 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25897 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25901 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25908 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25916 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25920 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25927 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25939 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25943 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25952 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25960 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25966 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25977 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_25985 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25989 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_25996 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26004 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26008 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26017 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26025 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26031 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26042 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26050 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26054 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26061 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26069 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26073 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26082 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26090 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26096 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26107 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26115 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26119 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26126 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26134 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26138 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26145 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26153 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26157 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26164 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26176 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26180 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26189 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26197 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26203 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26214 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26222 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26226 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26233 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26241 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26245 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26254 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26262 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26268 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26279 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26287 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26291 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26298 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26306 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26310 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26319 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26327 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26333 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26344 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26352 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26356 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26363 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26371 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26375 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26382 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26390 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26394 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26401 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26413 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26417 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26426 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26434 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26440 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26451 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26459 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26463 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26470 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26478 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26482 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26491 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26499 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26505 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26516 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26524 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26528 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26535 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26543 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26547 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26554 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26562 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26566 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26575 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26583 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26589 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26600 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26608 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26612 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26619 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26627 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26631 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26638 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26650 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26654 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26663 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26671 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26677 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26688 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26696 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26700 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26707 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26715 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26719 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26728 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26736 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26742 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26753 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26761 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26765 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26772 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26780 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26784 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26791 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26799 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26803 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26812 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26820 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26826 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26837 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26845 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26849 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26856 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26864 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26868 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26875 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26887 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26891 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26900 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26908 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26914 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26925 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26933 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26937 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26944 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26952 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26956 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26965 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26973 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26979 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_26990 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_26998 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27002 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27009 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27017 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27021 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27030 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27038 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27044 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27055 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27063 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27067 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27074 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27082 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27086 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27093 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27101 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27105 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27112 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27124 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27128 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27137 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27145 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27151 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27162 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27170 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27174 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27181 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27189 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27193 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27200 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27208 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27212 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27221 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27229 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27235 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27246 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27254 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27258 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27265 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27273 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27277 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27284 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27296 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27300 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27309 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27317 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27323 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27334 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27342 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27346 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27353 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27361 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27365 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27372 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27380 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27384 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27393 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27401 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27407 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27418 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27426 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27430 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27437 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27445 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27449 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27456 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27468 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27472 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27481 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27489 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27495 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27506 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27514 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27518 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27525 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27533 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27537 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27546 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27554 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27560 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27571 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27579 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27583 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27590 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27598 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27602 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27609 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27617 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27621 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27628 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27640 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27644 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27651 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27659 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27663 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27672 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27680 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27686 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27697 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27705 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27709 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27716 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27724 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27728 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27735 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27747 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27751 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27758 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27766 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27770 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27779 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27787 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27793 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27804 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27812 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27816 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27823 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27831 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27835 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27842 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27854 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27858 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27865 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27873 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27877 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27886 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27894 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27900 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27911 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27919 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27923 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27930 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27938 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27942 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27949 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27961 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27965 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27972 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_27980 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27984 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_27993 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28001 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28007 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28018 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28026 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28030 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28037 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28045 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28049 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28056 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28068 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28072 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28079 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28087 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28091 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28100 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28108 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28114 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28125 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28133 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28137 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28144 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28152 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28156 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28163 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28175 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28179 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28186 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28194 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28198 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28207 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28215 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28221 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28232 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28240 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28244 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28251 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28259 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28263 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28270 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28282 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28286 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28293 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28301 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28305 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28314 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28322 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28328 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28339 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28347 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28351 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28358 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28366 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28370 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28377 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28389 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28393 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28402 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28410 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28416 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28427 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28435 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28439 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28446 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28454 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28458 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28465 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28473 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28477 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28484 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28496 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28500 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28509 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28517 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28523 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28534 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28542 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28546 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28553 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28561 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28565 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28572 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28580 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28584 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28591 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28603 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28607 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28614 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28622 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28626 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28635 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28643 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28649 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28660 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28668 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28672 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28679 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28687 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28691 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28698 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28710 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28714 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28721 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28729 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28733 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28742 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28750 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28756 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28767 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28775 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28779 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28786 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28794 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28798 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28805 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28817 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28821 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28830 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28838 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28844 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28855 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28863 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28867 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28874 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28882 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28886 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28893 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28901 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28905 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28912 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28924 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28928 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28935 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28943 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28947 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28956 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28964 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28970 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28981 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_28989 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_28993 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29000 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29008 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29012 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29019 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29031 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29035 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29044 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29052 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29058 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29069 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29077 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29081 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29088 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29096 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29100 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29107 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29115 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29119 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29126 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29138 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29142 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29151 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29159 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29165 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29176 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29184 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29188 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29195 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29203 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29207 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29214 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29222 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29226 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29233 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29245 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29249 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29256 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29264 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29268 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29277 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29285 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29291 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29302 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29310 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29314 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29321 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29329 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29333 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29340 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29352 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29356 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29363 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29371 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29375 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29384 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29392 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29398 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29409 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29417 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29421 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29428 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29436 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29440 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29447 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29459 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29463 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29472 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29480 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29486 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29497 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29505 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29509 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29516 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29524 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29528 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29535 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29543 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29547 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29554 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29566 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29570 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29579 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29587 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29593 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29604 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29612 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29616 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29623 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29631 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29635 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29642 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29650 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29654 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29661 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29673 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29677 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29684 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29692 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29696 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29705 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29713 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29719 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29730 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29738 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29742 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29749 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29757 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29761 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29768 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29780 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29784 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29793 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29801 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29807 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29818 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29826 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29830 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29837 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29845 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29849 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29856 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29864 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29868 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29875 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29887 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29891 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29900 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29908 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29914 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29925 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29933 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29937 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29944 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29952 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29956 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29963 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29971 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29975 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29982 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_29994 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_29998 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30007 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30015 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30021 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30032 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30040 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30044 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30051 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30059 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30063 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30070 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30078 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30082 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30089 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30101 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30105 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30114 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30122 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30128 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30139 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30147 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30151 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30158 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30166 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30170 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30177 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30185 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30189 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30196 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30208 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30212 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30221 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30229 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30235 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30246 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30254 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30258 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30265 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30273 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30277 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30284 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30292 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30296 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30303 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30315 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30321 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30328 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30336 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30344 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30351 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30359 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30363 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30372 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30380 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30384 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30395 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30403 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30407 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30414 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30422 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30426 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30433 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30445 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30449 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30456 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30464 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30468 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30475 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30487 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30491 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30500 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30508 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30514 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30525 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30533 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30537 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30544 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30552 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30556 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30563 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30571 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30575 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30582 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30594 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30598 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30607 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30615 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30621 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30632 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30640 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30644 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30651 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30659 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30663 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30670 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30678 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30682 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30689 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30701 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30705 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30714 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30722 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30726 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30735 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30743 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30747 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30758 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30766 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30770 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30777 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30785 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30789 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30796 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30808 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30812 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30819 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30827 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30831 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30838 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30850 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30856 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30863 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30871 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30875 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30884 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30892 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30896 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30903 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30911 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30915 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30922 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30934 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30938 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30945 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30953 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30959 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30970 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30978 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30982 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_30989 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_30997 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31001 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31008 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31020 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31024 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31031 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31039 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31043 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31050 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31062 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31068 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31075 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31083 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31089 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31096 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31104 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31108 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31117 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31125 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31133 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31140 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31148 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31152 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31159 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31167 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31171 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31178 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31190 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31194 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31201 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31209 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31213 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31220 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31232 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31236 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31243 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31251 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31255 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31262 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31274 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31280 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31287 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31295 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31301 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31312 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31320 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31324 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31331 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31339 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31343 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31350 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31358 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31362 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31369 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31381 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31385 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31392 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31400 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31404 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31411 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31423 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31427 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31434 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31442 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31446 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31453 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31465 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31471 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31478 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31486 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31490 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31497 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31505 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31509 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31516 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31528 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31532 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31539 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31547 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31551 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31558 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31570 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31574 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31583 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31591 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31595 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31602 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31610 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31614 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31623 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31631 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31635 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31642 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31654 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31660 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31671 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31679 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31683 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31690 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31698 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31702 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31709 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31717 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31721 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31728 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31740 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31744 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31751 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31759 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31763 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31770 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31782 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31786 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31793 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31801 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31805 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31812 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31824 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31828 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31835 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31843 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31849 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31856 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31864 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31872 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31879 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31887 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31891 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31898 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31910 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31914 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31921 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31929 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31933 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31940 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31948 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31956 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31963 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31975 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31979 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31986 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_31994 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_31998 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32005 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32017 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32021 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32028 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32036 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32040 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32047 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32059 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32063 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32070 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32078 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32082 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32089 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32101 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32105 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32112 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32120 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32124 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32131 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32143 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32147 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32154 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32162 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32166 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32173 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32185 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32189 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32196 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32204 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32208 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32215 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32227 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32231 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32238 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32246 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32250 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32257 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32269 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32273 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32280 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32288 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32292 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32299 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32311 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32315 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32322 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32330 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32334 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32341 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32353 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32357 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32364 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32372 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32376 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32383 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32395 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32399 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32406 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32414 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32418 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32425 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32437 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32441 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32448 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32456 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32460 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32467 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32479 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32483 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32490 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32498 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32502 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32509 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32521 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32525 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32532 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32540 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32544 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32551 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32563 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32567 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32574 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32582 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32586 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32593 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32605 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32609 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32616 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32624 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32628 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32635 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32647 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32651 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32658 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32666 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32670 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32677 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32689 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32693 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32700 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32708 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32712 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32719 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32731 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32735 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32742 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32750 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32754 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32761 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32773 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32777 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32784 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32792 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32796 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32803 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32815 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32819 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32826 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32834 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32838 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32845 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32857 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32861 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32868 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32876 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32880 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32887 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32899 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32903 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32910 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32918 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32922 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32929 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32941 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32945 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32952 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32960 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32964 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32971 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_32983 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32987 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_32994 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33002 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33006 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33013 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33025 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33029 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33036 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33044 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33048 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33055 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33067 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33071 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33078 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33086 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33090 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33097 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33109 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33113 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33120 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33128 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33132 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33139 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33151 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33155 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33162 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33170 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33174 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33181 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33193 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33197 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33204 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33212 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33216 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33223 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33235 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33239 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33246 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33254 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33258 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33265 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33277 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33281 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33288 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33296 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33300 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33307 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33319 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33323 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33330 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33338 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33342 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33349 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33361 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33365 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33372 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33380 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33384 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33391 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33403 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33407 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33414 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33422 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33426 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33433 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33445 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33449 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33456 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33464 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33468 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33475 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33487 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33491 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33498 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33506 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33510 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33517 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33529 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33533 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33540 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33548 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33552 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33559 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33571 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33575 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33582 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33590 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33594 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33601 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33613 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33617 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33624 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33632 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33636 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33643 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33655 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33659 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33666 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33674 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33678 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33685 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33697 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33701 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33708 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33716 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33720 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33727 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33739 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33743 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33750 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33758 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33762 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33769 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33781 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33785 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33792 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33800 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33804 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33811 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33823 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33827 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33834 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33842 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33846 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33853 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33865 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33869 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33876 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33884 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33888 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33895 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33907 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33911 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33918 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33926 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33930 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33937 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33949 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33953 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33960 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33968 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33972 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33979 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_33991 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_33995 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34002 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34010 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34014 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34021 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34033 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34037 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34044 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34052 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34056 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34063 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34075 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34079 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34086 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34094 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34098 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34105 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34117 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34121 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34128 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34136 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34142 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34149 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34157 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34161 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34168 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34180 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34184 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34193 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34201 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34205 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34212 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34220 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34224 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34231 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34243 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34247 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34254 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34262 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34266 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34273 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34285 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34289 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34296 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34304 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34308 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34315 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34327 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34331 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34338 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34346 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34350 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34357 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34369 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34373 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34380 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34388 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34392 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34399 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34411 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34415 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34422 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34430 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34434 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34441 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34453 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34459 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34470 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34478 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34482 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34489 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34497 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34501 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34508 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34516 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34520 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34527 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34539 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34543 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34550 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34558 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34562 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34569 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34581 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34585 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34592 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34600 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34604 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34611 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34623 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34629 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34640 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34648 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34652 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34659 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34667 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34671 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34678 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34686 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34690 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34697 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34709 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34713 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34720 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34728 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34732 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34739 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34751 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34755 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34762 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34770 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34774 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34781 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34793 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34799 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34810 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34818 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34822 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34829 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34837 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34841 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34848 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34856 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34860 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34867 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34879 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34883 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34890 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34898 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34902 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34909 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34921 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34925 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34932 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34940 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34944 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34951 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34963 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34969 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34980 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_34988 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34992 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_34999 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35007 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35011 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35018 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35026 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35030 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35037 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35049 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35053 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35060 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35068 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35072 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35079 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35091 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35095 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35102 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35110 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35114 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35121 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35133 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35139 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35146 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35153 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35163 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35167 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35174 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35181 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35191 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35195 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35202 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35209 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35219 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35223 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35230 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35237 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35247 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35251 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35258 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35265 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35275 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35279 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35286 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35293 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35303 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35307 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35314 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35321 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35331 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35335 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35342 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35349 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35359 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35363 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35370 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35377 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35387 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35391 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35398 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35405 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35415 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35419 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35426 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35433 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35443 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35449 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35456 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35463 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35473 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35477 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35484 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35491 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35501 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35505 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35512 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35519 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35529 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35533 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35540 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35547 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35557 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35561 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35568 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35575 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35585 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35589 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35596 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35603 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35613 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35617 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35624 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35631 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35641 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35645 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35652 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35659 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35669 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35673 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35680 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35687 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35697 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35701 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35708 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35715 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35725 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35729 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35736 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35743 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35753 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35757 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35764 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35771 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35781 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35785 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35792 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35799 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35809 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35813 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35820 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35827 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35837 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35841 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35848 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35855 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35865 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35869 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35876 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35883 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35893 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35897 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35904 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35911 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35921 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35925 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35932 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35939 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35949 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35953 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35960 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35967 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_35977 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35981 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35988 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_35995 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36005 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36009 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36016 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36023 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36033 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36037 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36044 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36051 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36061 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36065 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36072 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36079 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36089 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36093 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36100 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36107 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36117 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36121 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36128 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36135 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36145 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36149 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36156 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36163 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36173 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36177 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36184 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36191 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36201 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36205 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36212 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36219 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36229 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36233 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36240 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36247 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36257 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36261 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36268 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36275 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36285 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36289 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36296 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36303 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36313 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36317 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36324 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36331 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36341 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36345 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36352 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36359 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36369 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36373 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36380 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36387 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36397 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36401 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36408 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36415 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36425 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36429 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36436 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36443 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36453 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36457 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36464 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36471 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36481 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36485 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36492 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36499 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36509 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36513 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36520 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36527 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36537 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36541 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36548 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36555 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36565 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36569 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36576 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36583 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36593 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36597 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36604 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36611 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36621 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36625 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36632 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36639 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36649 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36653 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36660 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36667 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36677 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36681 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36688 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36695 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36705 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36709 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36716 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36723 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36733 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36737 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36744 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36751 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36761 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36765 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36772 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36779 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36789 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36793 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36800 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36807 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36817 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36821 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36828 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36835 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36845 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36849 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36856 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36863 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36873 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36877 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36884 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36891 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36901 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36905 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36912 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36919 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36929 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36935 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36942 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36949 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36959 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36965 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36972 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36979 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_36989 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_36995 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37002 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37009 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37019 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37025 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37032 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37039 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37049 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37055 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37062 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37069 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37079 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37085 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37092 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37099 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37109 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37115 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37122 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37129 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37139 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37145 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37152 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37159 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37169 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37175 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37182 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37189 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37199 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37205 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37212 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37219 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37229 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37235 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37242 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37249 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37259 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37265 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37272 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37279 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37289 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37295 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37302 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37309 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37319 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37325 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37332 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37339 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37349 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37355 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37362 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37369 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37379 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37385 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37392 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37399 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37409 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37415 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37422 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37429 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37439 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37445 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37452 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37459 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37469 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37475 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37482 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37489 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37499 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37505 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37512 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37519 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37529 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37535 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37542 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37549 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37559 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37565 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37572 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37579 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37589 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37595 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37602 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37609 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37619 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37625 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37632 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37639 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37649 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37655 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37662 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37669 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37679 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37685 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37692 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37699 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37709 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37715 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37722 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37729 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37739 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37745 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37752 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37759 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37769 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37775 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37782 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37789 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37799 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37805 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37812 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37819 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37829 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37835 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37842 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37849 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37859 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37865 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37872 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37879 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37889 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37895 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37902 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37909 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37919 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37925 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37932 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37939 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37949 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37955 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37962 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37969 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_37979 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37985 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37992 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_37999 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38009 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38015 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38022 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38029 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38039 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38045 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38052 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38059 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38069 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38075 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38082 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38089 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38099 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38105 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38112 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38119 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38129 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38135 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38142 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38149 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38159 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38165 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38172 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38179 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38189 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38195 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38202 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38209 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38219 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38225 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38232 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38239 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38249 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38255 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38262 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38269 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38279 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38285 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38292 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38299 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38309 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38315 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38322 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38329 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38339 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38345 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38352 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38359 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38369 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38375 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38382 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38389 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38399 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38405 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38412 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38419 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38429 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38435 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38442 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38449 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38459 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38465 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38472 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38479 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38489 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38495 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38502 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38509 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38519 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38525 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38532 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38539 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38549 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38555 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38562 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38569 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38579 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38585 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38592 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38599 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38609 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38615 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38622 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38629 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38639 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38645 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38652 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38659 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38669 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38675 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38682 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38689 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38699 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38705 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38712 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38719 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38729 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38735 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38742 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38749 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38759 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38765 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38772 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38779 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38789 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38795 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38802 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38809 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38819 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38825 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38832 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38839 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38849 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38855 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38862 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38869 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38879 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38885 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38892 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38899 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38909 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38915 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38922 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38929 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38939 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38945 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38952 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38959 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38969 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38975 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38982 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_38989 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_38999 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39005 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39012 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39019 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39029 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39035 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39042 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39049 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39059 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39065 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39072 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39079 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39089 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39095 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39102 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39109 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39119 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39125 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39132 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39139 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39149 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39155 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39162 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39169 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39179 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39185 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39192 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39199 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39209 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39215 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39222 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39229 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39239 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39245 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39252 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39259 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39269 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39275 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39282 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39289 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39299 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39305 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39312 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39319 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39329 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39335 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39342 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39349 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39359 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39365 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39372 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39379 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39389 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39395 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39402 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39409 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39419 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39425 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39432 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39439 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39449 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39455 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39462 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39469 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39479 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39485 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39492 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39499 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39509 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39515 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39522 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39529 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39539 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39545 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39552 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39559 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39569 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39575 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39582 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39589 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39599 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39605 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39612 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39619 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39629 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39635 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39642 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39649 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39659 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39665 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39672 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39679 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39689 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39695 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39702 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39709 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39719 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39725 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39732 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39739 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39749 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39755 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39762 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39769 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39779 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39785 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39792 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39799 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39809 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39815 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39822 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39829 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39839 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39845 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39852 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39859 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39869 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39875 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39882 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39889 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39899 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39905 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39912 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39919 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39929 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39935 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39942 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39949 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39959 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39965 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39972 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39979 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_39989 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_39995 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40002 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40009 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40019 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40025 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40032 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40039 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40049 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40055 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40062 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40069 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40079 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40085 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40092 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40099 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40109 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40115 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40122 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40129 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40139 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40145 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40152 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40159 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40169 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40175 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40182 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40189 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40199 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40205 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40212 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40219 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40229 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40235 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40242 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40249 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40259 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40265 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40272 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40279 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40289 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40295 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40302 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40309 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40319 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40325 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40332 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40339 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40349 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40355 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40362 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40369 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40379 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40385 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40392 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40399 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40409 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40415 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40422 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40429 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40439 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40445 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40452 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40459 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40469 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40475 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40482 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40489 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40499 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40505 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40512 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40519 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40529 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40535 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40542 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40549 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40559 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40565 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40572 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40579 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40589 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40595 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40602 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40609 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40619 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40625 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40632 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40639 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40649 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40655 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40662 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40669 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40679 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40685 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40692 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40699 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40709 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40715 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40722 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40729 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40739 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40745 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40752 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40759 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40769 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40773 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40782 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40789 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40799 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40803 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40812 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40819 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40829 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40833 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40842 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40849 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40859 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40863 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40872 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40879 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40889 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40893 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40902 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40909 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40919 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40923 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40932 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40939 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40949 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40953 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40962 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40969 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_40979 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40983 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40992 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_40999 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41009 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41013 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41022 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41029 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41039 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41043 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41052 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41059 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41069 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41073 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41082 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41089 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41099 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41103 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41112 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41119 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41129 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41133 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41142 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41149 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41159 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41163 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41172 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41179 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41189 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41193 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41202 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41209 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41219 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41223 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41232 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41239 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41249 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41253 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41262 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41269 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41279 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41283 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41292 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41299 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41309 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41313 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41322 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41329 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41339 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41343 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41352 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41359 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41369 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41373 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41382 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41389 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41399 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41403 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41412 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41419 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41429 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41433 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41442 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41449 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41459 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41463 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41472 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41479 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41489 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41493 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41502 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41509 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41519 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41523 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41532 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41539 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41549 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41553 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41562 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41569 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41579 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41583 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41592 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41599 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41609 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41613 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41622 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41629 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41639 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41643 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41652 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41659 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41669 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41673 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41682 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41689 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41699 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41703 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41712 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41719 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41729 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41733 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41742 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41749 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41759 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41763 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41772 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41779 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41789 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41793 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41802 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41809 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41819 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41823 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41832 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41839 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41849 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41853 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41862 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41869 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41879 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41883 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41892 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41899 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41909 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41913 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41920 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41927 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41937 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41941 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41948 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41955 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41965 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41969 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41976 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41983 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_41993 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_41997 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42004 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42011 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42021 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42025 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42032 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42039 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42049 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42053 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42060 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42067 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42077 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42081 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42088 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42095 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42105 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42109 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42116 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42123 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42133 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42137 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42144 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42151 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42161 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42165 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42172 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42179 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42189 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42195 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42202 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42209 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42219 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42223 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42230 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42237 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42247 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42253 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42260 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42267 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42277 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42281 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42288 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42295 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42305 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42309 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42316 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42323 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42333 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42337 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42344 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42351 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42361 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42365 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42372 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42379 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42389 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42393 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42400 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42407 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42417 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42421 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42428 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42435 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42445 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42449 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42456 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42463 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42473 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42477 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42484 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42491 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42501 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42505 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42512 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42519 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42529 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42533 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42540 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42547 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42557 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42561 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42568 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42575 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42585 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42589 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42596 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42603 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42613 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42617 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42624 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42631 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42641 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42645 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42652 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42659 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42669 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42673 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42680 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42687 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42697 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42701 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42708 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42715 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42725 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42729 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42736 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42743 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42753 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42757 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42764 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42771 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42781 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42785 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42792 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42799 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42809 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42813 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42820 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42827 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42837 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42841 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42848 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42855 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42865 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42869 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42876 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42883 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42893 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42897 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42904 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42911 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42921 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42925 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42932 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42939 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42949 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42953 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42960 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42967 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_42977 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42981 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42988 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_42995 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43005 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43009 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43016 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43023 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43033 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43037 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43044 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43051 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43061 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43065 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43072 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43079 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43089 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43093 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43100 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43107 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43117 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43121 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43128 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43135 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43145 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43149 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43156 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43163 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43173 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43177 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43184 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43191 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43201 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43205 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43212 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43219 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43229 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43233 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43240 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43247 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43257 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43261 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43268 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43275 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43285 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43289 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43296 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43303 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43313 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43317 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43324 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43331 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43341 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43345 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43352 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43359 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43369 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43373 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43380 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43387 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43397 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43401 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43408 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43415 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43425 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43429 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43436 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43443 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43453 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43457 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43464 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43471 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43481 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43485 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43492 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43499 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43509 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43513 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43520 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43527 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43537 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43541 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43548 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43555 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43565 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43569 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43576 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43583 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43593 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43597 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43604 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43611 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43621 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43625 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43632 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43639 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43649 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43653 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43660 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43667 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43677 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43681 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43688 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43695 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43705 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43709 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43718 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43725 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43735 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43739 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43748 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43755 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43765 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43769 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43778 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43785 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43795 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43799 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43808 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43815 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43825 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43829 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43838 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43845 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43855 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43859 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43868 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43875 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43885 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43889 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43898 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43905 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43915 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43919 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43928 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43935 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43945 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43949 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43958 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43965 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_43975 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43979 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43988 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_43995 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44005 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44009 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44018 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44025 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44035 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44039 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44048 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44055 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44065 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44069 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44078 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44085 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44095 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44099 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44108 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44115 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44125 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44129 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44138 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44145 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44155 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44159 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44168 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44175 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44185 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44189 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44198 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44205 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44215 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44219 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44228 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44235 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44245 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44249 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44258 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44265 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44275 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44279 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44288 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44295 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44305 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44309 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44318 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44325 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44335 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44339 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44348 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44355 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44365 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44369 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44378 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44385 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44395 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44399 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44408 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44415 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44425 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44429 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44438 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44445 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44455 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44459 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44468 : std_logic_vector(2 downto 0);
  signal LPM_q_ivl_44475 : std_logic_vector(2 downto 0);
  signal LPM_d0_ivl_44485 : std_logic_vector(2 downto 0);
  
  component not_masked is
    port (
      a : in std_logic_vector(1 downto 0);
      b : out std_logic_vector(1 downto 0)
    );
  end component;
  
  component and_HPC2 is
    port (
      a : in std_logic_vector(2 downto 0);
      b : in std_logic_vector(2 downto 0);
      c : out std_logic_vector(2 downto 0);
      clk : in std_logic;
      r : in std_logic_vector(2 downto 0)
    );
  end component;
  
  component nor_HPC2 is
    port (
      a : in std_logic_vector(2 downto 0);
      b : in std_logic_vector(2 downto 0);
      c : out std_logic_vector(2 downto 0);
      clk : in std_logic;
      r : in std_logic_vector(2 downto 0)
    );
  end component;
  
  component xor_HPC2 is
    port (
      a : in std_logic_vector(2 downto 0);
      b : in std_logic_vector(2 downto 0);
      c : out std_logic_vector(2 downto 0)
    );
  end component;
  
  component xnor_HPC2 is
    port (
      a : in std_logic_vector(2 downto 0);
      b : in std_logic_vector(2 downto 0);
      c : out std_logic_vector(2 downto 0)
    );
  end component;
  
  component INV_X1 is
    port (
      A : in std_logic;
      ZN : out std_logic
    );
  end component;
  
  component XNOR2_X1 is
    port (
      A : in std_logic;
      B : in std_logic;
      ZN : out std_logic
    );
  end component;
  
  component NAND2_X1 is
    port (
      A1 : in std_logic;
      A2 : in std_logic;
      ZN : out std_logic
    );
  end component;
begin
  tmp_ivl_1 <= state_in_s1(241);
  tmp_ivl_3 <= state_in_s0(241);
  tmp_ivl_4 <= tmp_ivl_1 & tmp_ivl_3;
  LPM_q_ivl_7 <= tmp_ivl_9 & tmp_ivl_4;
  tmp_ivl_12 <= state_in_s1(305);
  tmp_ivl_14 <= state_in_s0(305);
  tmp_ivl_15 <= tmp_ivl_12 & tmp_ivl_14;
  LPM_q_ivl_18 <= tmp_ivl_20 & tmp_ivl_15;
  new_AGEMA_signal_2338 <= tmp_ivl_24(1);
  tmp_ivl_22 <= tmp_ivl_24(0);
  tmp_ivl_24 <= LPM_d0_ivl_28(0 + 1 downto 0);
  tmp_ivl_30 <= state_in_s1(304);
  tmp_ivl_32 <= state_in_s0(304);
  tmp_ivl_33 <= tmp_ivl_30 & tmp_ivl_32;
  LPM_q_ivl_36 <= tmp_ivl_38 & tmp_ivl_33;
  tmp_ivl_41 <= state_in_s1(240);
  tmp_ivl_43 <= state_in_s0(240);
  tmp_ivl_44 <= tmp_ivl_41 & tmp_ivl_43;
  LPM_q_ivl_47 <= tmp_ivl_49 & tmp_ivl_44;
  new_AGEMA_signal_2341 <= tmp_ivl_53(1);
  tmp_ivl_51 <= tmp_ivl_53(0);
  tmp_ivl_53 <= LPM_d0_ivl_57(0 + 1 downto 0);
  tmp_ivl_59 <= state_in_s1(255);
  tmp_ivl_61 <= state_in_s0(255);
  tmp_ivl_62 <= tmp_ivl_59 & tmp_ivl_61;
  LPM_q_ivl_65 <= tmp_ivl_67 & tmp_ivl_62;
  tmp_ivl_70 <= state_in_s1(319);
  tmp_ivl_72 <= state_in_s0(319);
  tmp_ivl_73 <= tmp_ivl_70 & tmp_ivl_72;
  LPM_q_ivl_76 <= tmp_ivl_78 & tmp_ivl_73;
  new_AGEMA_signal_2344 <= tmp_ivl_82(1);
  tmp_ivl_80 <= tmp_ivl_82(0);
  tmp_ivl_82 <= LPM_d0_ivl_86(0 + 1 downto 0);
  tmp_ivl_88 <= state_in_s1(254);
  tmp_ivl_90 <= state_in_s0(254);
  tmp_ivl_91 <= tmp_ivl_88 & tmp_ivl_90;
  LPM_q_ivl_94 <= tmp_ivl_96 & tmp_ivl_91;
  tmp_ivl_99 <= state_in_s1(318);
  tmp_ivl_101 <= state_in_s0(318);
  tmp_ivl_102 <= tmp_ivl_99 & tmp_ivl_101;
  LPM_q_ivl_105 <= tmp_ivl_107 & tmp_ivl_102;
  new_AGEMA_signal_2347 <= tmp_ivl_111(1);
  tmp_ivl_109 <= tmp_ivl_111(0);
  tmp_ivl_111 <= LPM_d0_ivl_115(0 + 1 downto 0);
  tmp_ivl_117 <= state_in_s1(199);
  tmp_ivl_119 <= state_in_s0(199);
  tmp_ivl_120 <= tmp_ivl_117 & tmp_ivl_119;
  LPM_q_ivl_123 <= tmp_ivl_125 & tmp_ivl_120;
  tmp_ivl_128 <= state_in_s1(263);
  tmp_ivl_130 <= state_in_s0(263);
  tmp_ivl_131 <= tmp_ivl_128 & tmp_ivl_130;
  LPM_q_ivl_134 <= tmp_ivl_136 & tmp_ivl_131;
  new_AGEMA_signal_2350 <= tmp_ivl_140(1);
  tmp_ivl_138 <= tmp_ivl_140(0);
  tmp_ivl_140 <= LPM_d0_ivl_144(0 + 1 downto 0);
  tmp_ivl_146 <= state_in_s1(262);
  tmp_ivl_148 <= state_in_s0(262);
  tmp_ivl_149 <= tmp_ivl_146 & tmp_ivl_148;
  LPM_q_ivl_152 <= tmp_ivl_154 & tmp_ivl_149;
  tmp_ivl_157 <= state_in_s1(198);
  tmp_ivl_159 <= state_in_s0(198);
  tmp_ivl_160 <= tmp_ivl_157 & tmp_ivl_159;
  LPM_q_ivl_163 <= tmp_ivl_165 & tmp_ivl_160;
  new_AGEMA_signal_2353 <= tmp_ivl_169(1);
  tmp_ivl_167 <= tmp_ivl_169(0);
  tmp_ivl_169 <= LPM_d0_ivl_173(0 + 1 downto 0);
  tmp_ivl_175 <= state_in_s1(197);
  tmp_ivl_177 <= state_in_s0(197);
  tmp_ivl_178 <= tmp_ivl_175 & tmp_ivl_177;
  LPM_q_ivl_181 <= tmp_ivl_183 & tmp_ivl_178;
  tmp_ivl_186 <= state_in_s1(261);
  tmp_ivl_188 <= state_in_s0(261);
  tmp_ivl_189 <= tmp_ivl_186 & tmp_ivl_188;
  LPM_q_ivl_192 <= tmp_ivl_194 & tmp_ivl_189;
  new_AGEMA_signal_2356 <= tmp_ivl_198(1);
  tmp_ivl_196 <= tmp_ivl_198(0);
  tmp_ivl_198 <= LPM_d0_ivl_202(0 + 1 downto 0);
  tmp_ivl_204 <= state_in_s1(196);
  tmp_ivl_206 <= state_in_s0(196);
  tmp_ivl_207 <= tmp_ivl_204 & tmp_ivl_206;
  LPM_q_ivl_210 <= tmp_ivl_212 & tmp_ivl_207;
  tmp_ivl_215 <= state_in_s1(260);
  tmp_ivl_217 <= state_in_s0(260);
  tmp_ivl_218 <= tmp_ivl_215 & tmp_ivl_217;
  LPM_q_ivl_221 <= tmp_ivl_223 & tmp_ivl_218;
  new_AGEMA_signal_2359 <= tmp_ivl_227(1);
  tmp_ivl_225 <= tmp_ivl_227(0);
  tmp_ivl_227 <= LPM_d0_ivl_231(0 + 1 downto 0);
  tmp_ivl_233 <= state_in_s1(317);
  tmp_ivl_235 <= state_in_s0(317);
  tmp_ivl_236 <= tmp_ivl_233 & tmp_ivl_235;
  LPM_q_ivl_239 <= tmp_ivl_241 & tmp_ivl_236;
  tmp_ivl_244 <= state_in_s1(253);
  tmp_ivl_246 <= state_in_s0(253);
  tmp_ivl_247 <= tmp_ivl_244 & tmp_ivl_246;
  LPM_q_ivl_250 <= tmp_ivl_252 & tmp_ivl_247;
  new_AGEMA_signal_2362 <= tmp_ivl_256(1);
  tmp_ivl_254 <= tmp_ivl_256(0);
  tmp_ivl_256 <= LPM_d0_ivl_260(0 + 1 downto 0);
  tmp_ivl_262 <= state_in_s1(195);
  tmp_ivl_264 <= state_in_s0(195);
  tmp_ivl_265 <= tmp_ivl_262 & tmp_ivl_264;
  LPM_q_ivl_268 <= tmp_ivl_270 & tmp_ivl_265;
  tmp_ivl_273 <= state_in_s1(259);
  tmp_ivl_275 <= state_in_s0(259);
  tmp_ivl_276 <= tmp_ivl_273 & tmp_ivl_275;
  LPM_q_ivl_279 <= tmp_ivl_281 & tmp_ivl_276;
  new_AGEMA_signal_2365 <= tmp_ivl_285(1);
  tmp_ivl_283 <= tmp_ivl_285(0);
  tmp_ivl_285 <= LPM_d0_ivl_289(0 + 1 downto 0);
  tmp_ivl_291 <= state_in_s1(258);
  tmp_ivl_293 <= state_in_s0(258);
  tmp_ivl_294 <= tmp_ivl_291 & tmp_ivl_293;
  LPM_q_ivl_297 <= tmp_ivl_299 & tmp_ivl_294;
  tmp_ivl_302 <= state_in_s1(194);
  tmp_ivl_304 <= state_in_s0(194);
  tmp_ivl_305 <= tmp_ivl_302 & tmp_ivl_304;
  LPM_q_ivl_308 <= tmp_ivl_310 & tmp_ivl_305;
  new_AGEMA_signal_2368 <= tmp_ivl_314(1);
  tmp_ivl_312 <= tmp_ivl_314(0);
  tmp_ivl_314 <= LPM_d0_ivl_318(0 + 1 downto 0);
  tmp_ivl_320 <= state_in_s1(193);
  tmp_ivl_322 <= state_in_s0(193);
  tmp_ivl_323 <= tmp_ivl_320 & tmp_ivl_322;
  LPM_q_ivl_326 <= tmp_ivl_328 & tmp_ivl_323;
  tmp_ivl_331 <= state_in_s1(257);
  tmp_ivl_333 <= state_in_s0(257);
  tmp_ivl_334 <= tmp_ivl_331 & tmp_ivl_333;
  LPM_q_ivl_337 <= tmp_ivl_339 & tmp_ivl_334;
  new_AGEMA_signal_2371 <= tmp_ivl_343(1);
  tmp_ivl_341 <= tmp_ivl_343(0);
  tmp_ivl_343 <= LPM_d0_ivl_347(0 + 1 downto 0);
  tmp_ivl_349 <= state_in_s1(192);
  tmp_ivl_351 <= state_in_s0(192);
  tmp_ivl_352 <= tmp_ivl_349 & tmp_ivl_351;
  LPM_q_ivl_355 <= tmp_ivl_357 & tmp_ivl_352;
  tmp_ivl_360 <= state_in_s1(256);
  tmp_ivl_362 <= state_in_s0(256);
  tmp_ivl_363 <= tmp_ivl_360 & tmp_ivl_362;
  LPM_q_ivl_366 <= tmp_ivl_368 & tmp_ivl_363;
  new_AGEMA_signal_2374 <= tmp_ivl_372(1);
  tmp_ivl_370 <= tmp_ivl_372(0);
  tmp_ivl_372 <= LPM_d0_ivl_376(0 + 1 downto 0);
  tmp_ivl_378 <= state_in_s1(271);
  tmp_ivl_380 <= state_in_s0(271);
  tmp_ivl_381 <= tmp_ivl_378 & tmp_ivl_380;
  LPM_q_ivl_384 <= tmp_ivl_386 & tmp_ivl_381;
  tmp_ivl_389 <= state_in_s1(207);
  tmp_ivl_391 <= state_in_s0(207);
  tmp_ivl_392 <= tmp_ivl_389 & tmp_ivl_391;
  LPM_q_ivl_395 <= tmp_ivl_397 & tmp_ivl_392;
  new_AGEMA_signal_2377 <= tmp_ivl_401(1);
  tmp_ivl_399 <= tmp_ivl_401(0);
  tmp_ivl_401 <= LPM_d0_ivl_405(0 + 1 downto 0);
  tmp_ivl_407 <= state_in_s1(206);
  tmp_ivl_409 <= state_in_s0(206);
  tmp_ivl_410 <= tmp_ivl_407 & tmp_ivl_409;
  LPM_q_ivl_413 <= tmp_ivl_415 & tmp_ivl_410;
  tmp_ivl_418 <= state_in_s1(270);
  tmp_ivl_420 <= state_in_s0(270);
  tmp_ivl_421 <= tmp_ivl_418 & tmp_ivl_420;
  LPM_q_ivl_424 <= tmp_ivl_426 & tmp_ivl_421;
  new_AGEMA_signal_2380 <= tmp_ivl_430(1);
  tmp_ivl_428 <= tmp_ivl_430(0);
  tmp_ivl_430 <= LPM_d0_ivl_434(0 + 1 downto 0);
  tmp_ivl_436 <= state_in_s1(205);
  tmp_ivl_438 <= state_in_s0(205);
  tmp_ivl_439 <= tmp_ivl_436 & tmp_ivl_438;
  LPM_q_ivl_442 <= tmp_ivl_444 & tmp_ivl_439;
  tmp_ivl_447 <= state_in_s1(269);
  tmp_ivl_449 <= state_in_s0(269);
  tmp_ivl_450 <= tmp_ivl_447 & tmp_ivl_449;
  LPM_q_ivl_453 <= tmp_ivl_455 & tmp_ivl_450;
  new_AGEMA_signal_2383 <= tmp_ivl_459(1);
  tmp_ivl_457 <= tmp_ivl_459(0);
  tmp_ivl_459 <= LPM_d0_ivl_463(0 + 1 downto 0);
  tmp_ivl_465 <= state_in_s1(268);
  tmp_ivl_467 <= state_in_s0(268);
  tmp_ivl_468 <= tmp_ivl_465 & tmp_ivl_467;
  LPM_q_ivl_471 <= tmp_ivl_473 & tmp_ivl_468;
  tmp_ivl_476 <= state_in_s1(204);
  tmp_ivl_478 <= state_in_s0(204);
  tmp_ivl_479 <= tmp_ivl_476 & tmp_ivl_478;
  LPM_q_ivl_482 <= tmp_ivl_484 & tmp_ivl_479;
  new_AGEMA_signal_2386 <= tmp_ivl_488(1);
  tmp_ivl_486 <= tmp_ivl_488(0);
  tmp_ivl_488 <= LPM_d0_ivl_492(0 + 1 downto 0);
  tmp_ivl_494 <= state_in_s1(267);
  tmp_ivl_496 <= state_in_s0(267);
  tmp_ivl_497 <= tmp_ivl_494 & tmp_ivl_496;
  LPM_q_ivl_500 <= tmp_ivl_502 & tmp_ivl_497;
  tmp_ivl_505 <= state_in_s1(203);
  tmp_ivl_507 <= state_in_s0(203);
  tmp_ivl_508 <= tmp_ivl_505 & tmp_ivl_507;
  LPM_q_ivl_511 <= tmp_ivl_513 & tmp_ivl_508;
  new_AGEMA_signal_2389 <= tmp_ivl_517(1);
  tmp_ivl_515 <= tmp_ivl_517(0);
  tmp_ivl_517 <= LPM_d0_ivl_521(0 + 1 downto 0);
  tmp_ivl_523 <= state_in_s1(202);
  tmp_ivl_525 <= state_in_s0(202);
  tmp_ivl_526 <= tmp_ivl_523 & tmp_ivl_525;
  LPM_q_ivl_529 <= tmp_ivl_531 & tmp_ivl_526;
  tmp_ivl_534 <= state_in_s1(266);
  tmp_ivl_536 <= state_in_s0(266);
  tmp_ivl_537 <= tmp_ivl_534 & tmp_ivl_536;
  LPM_q_ivl_540 <= tmp_ivl_542 & tmp_ivl_537;
  new_AGEMA_signal_2392 <= tmp_ivl_546(1);
  tmp_ivl_544 <= tmp_ivl_546(0);
  tmp_ivl_546 <= LPM_d0_ivl_550(0 + 1 downto 0);
  tmp_ivl_552 <= state_in_s1(316);
  tmp_ivl_554 <= state_in_s0(316);
  tmp_ivl_555 <= tmp_ivl_552 & tmp_ivl_554;
  LPM_q_ivl_558 <= tmp_ivl_560 & tmp_ivl_555;
  tmp_ivl_563 <= state_in_s1(252);
  tmp_ivl_565 <= state_in_s0(252);
  tmp_ivl_566 <= tmp_ivl_563 & tmp_ivl_565;
  LPM_q_ivl_569 <= tmp_ivl_571 & tmp_ivl_566;
  new_AGEMA_signal_2395 <= tmp_ivl_575(1);
  tmp_ivl_573 <= tmp_ivl_575(0);
  tmp_ivl_575 <= LPM_d0_ivl_579(0 + 1 downto 0);
  tmp_ivl_581 <= state_in_s1(201);
  tmp_ivl_583 <= state_in_s0(201);
  tmp_ivl_584 <= tmp_ivl_581 & tmp_ivl_583;
  LPM_q_ivl_587 <= tmp_ivl_589 & tmp_ivl_584;
  tmp_ivl_592 <= state_in_s1(265);
  tmp_ivl_594 <= state_in_s0(265);
  tmp_ivl_595 <= tmp_ivl_592 & tmp_ivl_594;
  LPM_q_ivl_598 <= tmp_ivl_600 & tmp_ivl_595;
  new_AGEMA_signal_2398 <= tmp_ivl_604(1);
  tmp_ivl_602 <= tmp_ivl_604(0);
  tmp_ivl_604 <= LPM_d0_ivl_608(0 + 1 downto 0);
  tmp_ivl_610 <= state_in_s1(264);
  tmp_ivl_612 <= state_in_s0(264);
  tmp_ivl_613 <= tmp_ivl_610 & tmp_ivl_612;
  LPM_q_ivl_616 <= tmp_ivl_618 & tmp_ivl_613;
  tmp_ivl_621 <= state_in_s1(200);
  tmp_ivl_623 <= state_in_s0(200);
  tmp_ivl_624 <= tmp_ivl_621 & tmp_ivl_623;
  LPM_q_ivl_627 <= tmp_ivl_629 & tmp_ivl_624;
  new_AGEMA_signal_2401 <= tmp_ivl_633(1);
  tmp_ivl_631 <= tmp_ivl_633(0);
  tmp_ivl_633 <= LPM_d0_ivl_637(0 + 1 downto 0);
  tmp_ivl_639 <= state_in_s1(279);
  tmp_ivl_641 <= state_in_s0(279);
  tmp_ivl_642 <= tmp_ivl_639 & tmp_ivl_641;
  LPM_q_ivl_645 <= tmp_ivl_647 & tmp_ivl_642;
  tmp_ivl_650 <= state_in_s1(215);
  tmp_ivl_652 <= state_in_s0(215);
  tmp_ivl_653 <= tmp_ivl_650 & tmp_ivl_652;
  LPM_q_ivl_656 <= tmp_ivl_658 & tmp_ivl_653;
  new_AGEMA_signal_2404 <= tmp_ivl_662(1);
  tmp_ivl_660 <= tmp_ivl_662(0);
  tmp_ivl_662 <= LPM_d0_ivl_666(0 + 1 downto 0);
  tmp_ivl_668 <= state_in_s1(278);
  tmp_ivl_670 <= state_in_s0(278);
  tmp_ivl_671 <= tmp_ivl_668 & tmp_ivl_670;
  LPM_q_ivl_674 <= tmp_ivl_676 & tmp_ivl_671;
  tmp_ivl_679 <= state_in_s1(214);
  tmp_ivl_681 <= state_in_s0(214);
  tmp_ivl_682 <= tmp_ivl_679 & tmp_ivl_681;
  LPM_q_ivl_685 <= tmp_ivl_687 & tmp_ivl_682;
  new_AGEMA_signal_2407 <= tmp_ivl_691(1);
  tmp_ivl_689 <= tmp_ivl_691(0);
  tmp_ivl_691 <= LPM_d0_ivl_695(0 + 1 downto 0);
  tmp_ivl_697 <= state_in_s1(277);
  tmp_ivl_699 <= state_in_s0(277);
  tmp_ivl_700 <= tmp_ivl_697 & tmp_ivl_699;
  LPM_q_ivl_703 <= tmp_ivl_705 & tmp_ivl_700;
  tmp_ivl_708 <= state_in_s1(213);
  tmp_ivl_710 <= state_in_s0(213);
  tmp_ivl_711 <= tmp_ivl_708 & tmp_ivl_710;
  LPM_q_ivl_714 <= tmp_ivl_716 & tmp_ivl_711;
  new_AGEMA_signal_2410 <= tmp_ivl_720(1);
  tmp_ivl_718 <= tmp_ivl_720(0);
  tmp_ivl_720 <= LPM_d0_ivl_724(0 + 1 downto 0);
  tmp_ivl_726 <= state_in_s1(276);
  tmp_ivl_728 <= state_in_s0(276);
  tmp_ivl_729 <= tmp_ivl_726 & tmp_ivl_728;
  LPM_q_ivl_732 <= tmp_ivl_734 & tmp_ivl_729;
  tmp_ivl_737 <= state_in_s1(212);
  tmp_ivl_739 <= state_in_s0(212);
  tmp_ivl_740 <= tmp_ivl_737 & tmp_ivl_739;
  LPM_q_ivl_743 <= tmp_ivl_745 & tmp_ivl_740;
  new_AGEMA_signal_2413 <= tmp_ivl_749(1);
  tmp_ivl_747 <= tmp_ivl_749(0);
  tmp_ivl_749 <= LPM_d0_ivl_753(0 + 1 downto 0);
  tmp_ivl_755 <= state_in_s1(275);
  tmp_ivl_757 <= state_in_s0(275);
  tmp_ivl_758 <= tmp_ivl_755 & tmp_ivl_757;
  LPM_q_ivl_761 <= tmp_ivl_763 & tmp_ivl_758;
  tmp_ivl_766 <= state_in_s1(211);
  tmp_ivl_768 <= state_in_s0(211);
  tmp_ivl_769 <= tmp_ivl_766 & tmp_ivl_768;
  LPM_q_ivl_772 <= tmp_ivl_774 & tmp_ivl_769;
  new_AGEMA_signal_2416 <= tmp_ivl_778(1);
  tmp_ivl_776 <= tmp_ivl_778(0);
  tmp_ivl_778 <= LPM_d0_ivl_782(0 + 1 downto 0);
  tmp_ivl_784 <= state_in_s1(274);
  tmp_ivl_786 <= state_in_s0(274);
  tmp_ivl_787 <= tmp_ivl_784 & tmp_ivl_786;
  LPM_q_ivl_790 <= tmp_ivl_792 & tmp_ivl_787;
  tmp_ivl_795 <= state_in_s1(210);
  tmp_ivl_797 <= state_in_s0(210);
  tmp_ivl_798 <= tmp_ivl_795 & tmp_ivl_797;
  LPM_q_ivl_801 <= tmp_ivl_803 & tmp_ivl_798;
  new_AGEMA_signal_2419 <= tmp_ivl_807(1);
  tmp_ivl_805 <= tmp_ivl_807(0);
  tmp_ivl_807 <= LPM_d0_ivl_811(0 + 1 downto 0);
  tmp_ivl_813 <= state_in_s1(273);
  tmp_ivl_815 <= state_in_s0(273);
  tmp_ivl_816 <= tmp_ivl_813 & tmp_ivl_815;
  LPM_q_ivl_819 <= tmp_ivl_821 & tmp_ivl_816;
  tmp_ivl_824 <= state_in_s1(209);
  tmp_ivl_826 <= state_in_s0(209);
  tmp_ivl_827 <= tmp_ivl_824 & tmp_ivl_826;
  LPM_q_ivl_830 <= tmp_ivl_832 & tmp_ivl_827;
  new_AGEMA_signal_2422 <= tmp_ivl_836(1);
  tmp_ivl_834 <= tmp_ivl_836(0);
  tmp_ivl_836 <= LPM_d0_ivl_840(0 + 1 downto 0);
  tmp_ivl_842 <= state_in_s1(272);
  tmp_ivl_844 <= state_in_s0(272);
  tmp_ivl_845 <= tmp_ivl_842 & tmp_ivl_844;
  LPM_q_ivl_848 <= tmp_ivl_850 & tmp_ivl_845;
  tmp_ivl_853 <= state_in_s1(208);
  tmp_ivl_855 <= state_in_s0(208);
  tmp_ivl_856 <= tmp_ivl_853 & tmp_ivl_855;
  LPM_q_ivl_859 <= tmp_ivl_861 & tmp_ivl_856;
  new_AGEMA_signal_2425 <= tmp_ivl_865(1);
  tmp_ivl_863 <= tmp_ivl_865(0);
  tmp_ivl_865 <= LPM_d0_ivl_869(0 + 1 downto 0);
  tmp_ivl_871 <= state_in_s1(251);
  tmp_ivl_873 <= state_in_s0(251);
  tmp_ivl_874 <= tmp_ivl_871 & tmp_ivl_873;
  LPM_q_ivl_877 <= tmp_ivl_879 & tmp_ivl_874;
  tmp_ivl_882 <= state_in_s1(315);
  tmp_ivl_884 <= state_in_s0(315);
  tmp_ivl_885 <= tmp_ivl_882 & tmp_ivl_884;
  LPM_q_ivl_888 <= tmp_ivl_890 & tmp_ivl_885;
  new_AGEMA_signal_2428 <= tmp_ivl_894(1);
  tmp_ivl_892 <= tmp_ivl_894(0);
  tmp_ivl_894 <= LPM_d0_ivl_898(0 + 1 downto 0);
  tmp_ivl_900 <= state_in_s1(287);
  tmp_ivl_902 <= state_in_s0(287);
  tmp_ivl_903 <= tmp_ivl_900 & tmp_ivl_902;
  LPM_q_ivl_906 <= tmp_ivl_908 & tmp_ivl_903;
  tmp_ivl_911 <= state_in_s1(223);
  tmp_ivl_913 <= state_in_s0(223);
  tmp_ivl_914 <= tmp_ivl_911 & tmp_ivl_913;
  LPM_q_ivl_917 <= tmp_ivl_919 & tmp_ivl_914;
  new_AGEMA_signal_2431 <= tmp_ivl_923(1);
  tmp_ivl_921 <= tmp_ivl_923(0);
  tmp_ivl_923 <= LPM_d0_ivl_927(0 + 1 downto 0);
  tmp_ivl_929 <= state_in_s1(286);
  tmp_ivl_931 <= state_in_s0(286);
  tmp_ivl_932 <= tmp_ivl_929 & tmp_ivl_931;
  LPM_q_ivl_935 <= tmp_ivl_937 & tmp_ivl_932;
  tmp_ivl_940 <= state_in_s1(222);
  tmp_ivl_942 <= state_in_s0(222);
  tmp_ivl_943 <= tmp_ivl_940 & tmp_ivl_942;
  LPM_q_ivl_946 <= tmp_ivl_948 & tmp_ivl_943;
  new_AGEMA_signal_2434 <= tmp_ivl_952(1);
  tmp_ivl_950 <= tmp_ivl_952(0);
  tmp_ivl_952 <= LPM_d0_ivl_956(0 + 1 downto 0);
  tmp_ivl_958 <= state_in_s1(285);
  tmp_ivl_960 <= state_in_s0(285);
  tmp_ivl_961 <= tmp_ivl_958 & tmp_ivl_960;
  LPM_q_ivl_964 <= tmp_ivl_966 & tmp_ivl_961;
  tmp_ivl_969 <= state_in_s1(221);
  tmp_ivl_971 <= state_in_s0(221);
  tmp_ivl_972 <= tmp_ivl_969 & tmp_ivl_971;
  LPM_q_ivl_975 <= tmp_ivl_977 & tmp_ivl_972;
  new_AGEMA_signal_2437 <= tmp_ivl_981(1);
  tmp_ivl_979 <= tmp_ivl_981(0);
  tmp_ivl_981 <= LPM_d0_ivl_985(0 + 1 downto 0);
  tmp_ivl_987 <= state_in_s1(284);
  tmp_ivl_989 <= state_in_s0(284);
  tmp_ivl_990 <= tmp_ivl_987 & tmp_ivl_989;
  LPM_q_ivl_993 <= tmp_ivl_995 & tmp_ivl_990;
  tmp_ivl_998 <= state_in_s1(220);
  tmp_ivl_1000 <= state_in_s0(220);
  tmp_ivl_1001 <= tmp_ivl_998 & tmp_ivl_1000;
  LPM_q_ivl_1004 <= tmp_ivl_1006 & tmp_ivl_1001;
  new_AGEMA_signal_2440 <= tmp_ivl_1010(1);
  tmp_ivl_1008 <= tmp_ivl_1010(0);
  tmp_ivl_1010 <= LPM_d0_ivl_1014(0 + 1 downto 0);
  tmp_ivl_1016 <= state_in_s1(283);
  tmp_ivl_1018 <= state_in_s0(283);
  tmp_ivl_1019 <= tmp_ivl_1016 & tmp_ivl_1018;
  LPM_q_ivl_1022 <= tmp_ivl_1024 & tmp_ivl_1019;
  tmp_ivl_1027 <= state_in_s1(219);
  tmp_ivl_1029 <= state_in_s0(219);
  tmp_ivl_1030 <= tmp_ivl_1027 & tmp_ivl_1029;
  LPM_q_ivl_1033 <= tmp_ivl_1035 & tmp_ivl_1030;
  new_AGEMA_signal_2443 <= tmp_ivl_1039(1);
  tmp_ivl_1037 <= tmp_ivl_1039(0);
  tmp_ivl_1039 <= LPM_d0_ivl_1043(0 + 1 downto 0);
  tmp_ivl_1045 <= state_in_s1(282);
  tmp_ivl_1047 <= state_in_s0(282);
  tmp_ivl_1048 <= tmp_ivl_1045 & tmp_ivl_1047;
  LPM_q_ivl_1051 <= tmp_ivl_1053 & tmp_ivl_1048;
  tmp_ivl_1056 <= state_in_s1(218);
  tmp_ivl_1058 <= state_in_s0(218);
  tmp_ivl_1059 <= tmp_ivl_1056 & tmp_ivl_1058;
  LPM_q_ivl_1062 <= tmp_ivl_1064 & tmp_ivl_1059;
  new_AGEMA_signal_2446 <= tmp_ivl_1068(1);
  tmp_ivl_1066 <= tmp_ivl_1068(0);
  tmp_ivl_1068 <= LPM_d0_ivl_1072(0 + 1 downto 0);
  tmp_ivl_1074 <= state_in_s1(281);
  tmp_ivl_1076 <= state_in_s0(281);
  tmp_ivl_1077 <= tmp_ivl_1074 & tmp_ivl_1076;
  LPM_q_ivl_1080 <= tmp_ivl_1082 & tmp_ivl_1077;
  tmp_ivl_1085 <= state_in_s1(217);
  tmp_ivl_1087 <= state_in_s0(217);
  tmp_ivl_1088 <= tmp_ivl_1085 & tmp_ivl_1087;
  LPM_q_ivl_1091 <= tmp_ivl_1093 & tmp_ivl_1088;
  new_AGEMA_signal_2449 <= tmp_ivl_1097(1);
  tmp_ivl_1095 <= tmp_ivl_1097(0);
  tmp_ivl_1097 <= LPM_d0_ivl_1101(0 + 1 downto 0);
  tmp_ivl_1103 <= state_in_s1(280);
  tmp_ivl_1105 <= state_in_s0(280);
  tmp_ivl_1106 <= tmp_ivl_1103 & tmp_ivl_1105;
  LPM_q_ivl_1109 <= tmp_ivl_1111 & tmp_ivl_1106;
  tmp_ivl_1114 <= state_in_s1(216);
  tmp_ivl_1116 <= state_in_s0(216);
  tmp_ivl_1117 <= tmp_ivl_1114 & tmp_ivl_1116;
  LPM_q_ivl_1120 <= tmp_ivl_1122 & tmp_ivl_1117;
  new_AGEMA_signal_2452 <= tmp_ivl_1126(1);
  tmp_ivl_1124 <= tmp_ivl_1126(0);
  tmp_ivl_1126 <= LPM_d0_ivl_1130(0 + 1 downto 0);
  tmp_ivl_1132 <= state_in_s1(295);
  tmp_ivl_1134 <= state_in_s0(295);
  tmp_ivl_1135 <= tmp_ivl_1132 & tmp_ivl_1134;
  LPM_q_ivl_1138 <= tmp_ivl_1140 & tmp_ivl_1135;
  tmp_ivl_1143 <= state_in_s1(231);
  tmp_ivl_1145 <= state_in_s0(231);
  tmp_ivl_1146 <= tmp_ivl_1143 & tmp_ivl_1145;
  LPM_q_ivl_1149 <= tmp_ivl_1151 & tmp_ivl_1146;
  new_AGEMA_signal_2455 <= tmp_ivl_1155(1);
  tmp_ivl_1153 <= tmp_ivl_1155(0);
  tmp_ivl_1155 <= LPM_d0_ivl_1159(0 + 1 downto 0);
  tmp_ivl_1161 <= state_in_s1(294);
  tmp_ivl_1163 <= state_in_s0(294);
  tmp_ivl_1164 <= tmp_ivl_1161 & tmp_ivl_1163;
  LPM_q_ivl_1167 <= tmp_ivl_1169 & tmp_ivl_1164;
  tmp_ivl_1172 <= state_in_s1(230);
  tmp_ivl_1174 <= state_in_s0(230);
  tmp_ivl_1175 <= tmp_ivl_1172 & tmp_ivl_1174;
  LPM_q_ivl_1178 <= tmp_ivl_1180 & tmp_ivl_1175;
  new_AGEMA_signal_2458 <= tmp_ivl_1184(1);
  tmp_ivl_1182 <= tmp_ivl_1184(0);
  tmp_ivl_1184 <= LPM_d0_ivl_1188(0 + 1 downto 0);
  tmp_ivl_1190 <= state_in_s1(250);
  tmp_ivl_1192 <= state_in_s0(250);
  tmp_ivl_1193 <= tmp_ivl_1190 & tmp_ivl_1192;
  LPM_q_ivl_1196 <= tmp_ivl_1198 & tmp_ivl_1193;
  tmp_ivl_1201 <= state_in_s1(314);
  tmp_ivl_1203 <= state_in_s0(314);
  tmp_ivl_1204 <= tmp_ivl_1201 & tmp_ivl_1203;
  LPM_q_ivl_1207 <= tmp_ivl_1209 & tmp_ivl_1204;
  new_AGEMA_signal_2461 <= tmp_ivl_1213(1);
  tmp_ivl_1211 <= tmp_ivl_1213(0);
  tmp_ivl_1213 <= LPM_d0_ivl_1217(0 + 1 downto 0);
  tmp_ivl_1219 <= state_in_s1(293);
  tmp_ivl_1221 <= state_in_s0(293);
  tmp_ivl_1222 <= tmp_ivl_1219 & tmp_ivl_1221;
  LPM_q_ivl_1225 <= tmp_ivl_1227 & tmp_ivl_1222;
  tmp_ivl_1230 <= state_in_s1(229);
  tmp_ivl_1232 <= state_in_s0(229);
  tmp_ivl_1233 <= tmp_ivl_1230 & tmp_ivl_1232;
  LPM_q_ivl_1236 <= tmp_ivl_1238 & tmp_ivl_1233;
  new_AGEMA_signal_2464 <= tmp_ivl_1242(1);
  tmp_ivl_1240 <= tmp_ivl_1242(0);
  tmp_ivl_1242 <= LPM_d0_ivl_1246(0 + 1 downto 0);
  tmp_ivl_1248 <= state_in_s1(292);
  tmp_ivl_1250 <= state_in_s0(292);
  tmp_ivl_1251 <= tmp_ivl_1248 & tmp_ivl_1250;
  LPM_q_ivl_1254 <= tmp_ivl_1256 & tmp_ivl_1251;
  tmp_ivl_1259 <= state_in_s1(228);
  tmp_ivl_1261 <= state_in_s0(228);
  tmp_ivl_1262 <= tmp_ivl_1259 & tmp_ivl_1261;
  LPM_q_ivl_1265 <= tmp_ivl_1267 & tmp_ivl_1262;
  new_AGEMA_signal_2467 <= tmp_ivl_1271(1);
  tmp_ivl_1269 <= tmp_ivl_1271(0);
  tmp_ivl_1271 <= LPM_d0_ivl_1275(0 + 1 downto 0);
  tmp_ivl_1277 <= state_in_s1(291);
  tmp_ivl_1279 <= state_in_s0(291);
  tmp_ivl_1280 <= tmp_ivl_1277 & tmp_ivl_1279;
  LPM_q_ivl_1283 <= tmp_ivl_1285 & tmp_ivl_1280;
  tmp_ivl_1288 <= state_in_s1(227);
  tmp_ivl_1290 <= state_in_s0(227);
  tmp_ivl_1291 <= tmp_ivl_1288 & tmp_ivl_1290;
  LPM_q_ivl_1294 <= tmp_ivl_1296 & tmp_ivl_1291;
  new_AGEMA_signal_2470 <= tmp_ivl_1300(1);
  tmp_ivl_1298 <= tmp_ivl_1300(0);
  tmp_ivl_1300 <= LPM_d0_ivl_1304(0 + 1 downto 0);
  tmp_ivl_1306 <= state_in_s1(290);
  tmp_ivl_1308 <= state_in_s0(290);
  tmp_ivl_1309 <= tmp_ivl_1306 & tmp_ivl_1308;
  LPM_q_ivl_1312 <= tmp_ivl_1314 & tmp_ivl_1309;
  tmp_ivl_1317 <= state_in_s1(226);
  tmp_ivl_1319 <= state_in_s0(226);
  tmp_ivl_1320 <= tmp_ivl_1317 & tmp_ivl_1319;
  LPM_q_ivl_1323 <= tmp_ivl_1325 & tmp_ivl_1320;
  new_AGEMA_signal_2473 <= tmp_ivl_1329(1);
  tmp_ivl_1327 <= tmp_ivl_1329(0);
  tmp_ivl_1329 <= LPM_d0_ivl_1333(0 + 1 downto 0);
  tmp_ivl_1335 <= state_in_s1(289);
  tmp_ivl_1337 <= state_in_s0(289);
  tmp_ivl_1338 <= tmp_ivl_1335 & tmp_ivl_1337;
  LPM_q_ivl_1341 <= tmp_ivl_1343 & tmp_ivl_1338;
  tmp_ivl_1346 <= state_in_s1(225);
  tmp_ivl_1348 <= state_in_s0(225);
  tmp_ivl_1349 <= tmp_ivl_1346 & tmp_ivl_1348;
  LPM_q_ivl_1352 <= tmp_ivl_1354 & tmp_ivl_1349;
  new_AGEMA_signal_2476 <= tmp_ivl_1358(1);
  tmp_ivl_1356 <= tmp_ivl_1358(0);
  tmp_ivl_1358 <= LPM_d0_ivl_1362(0 + 1 downto 0);
  tmp_ivl_1364 <= state_in_s1(224);
  tmp_ivl_1366 <= state_in_s0(224);
  tmp_ivl_1367 <= tmp_ivl_1364 & tmp_ivl_1366;
  LPM_q_ivl_1370 <= tmp_ivl_1372 & tmp_ivl_1367;
  tmp_ivl_1375 <= state_in_s1(288);
  tmp_ivl_1377 <= state_in_s0(288);
  tmp_ivl_1378 <= tmp_ivl_1375 & tmp_ivl_1377;
  LPM_q_ivl_1381 <= tmp_ivl_1383 & tmp_ivl_1378;
  new_AGEMA_signal_2479 <= tmp_ivl_1387(1);
  tmp_ivl_1385 <= tmp_ivl_1387(0);
  tmp_ivl_1387 <= LPM_d0_ivl_1391(0 + 1 downto 0);
  tmp_ivl_1393 <= state_in_s1(239);
  tmp_ivl_1395 <= state_in_s0(239);
  tmp_ivl_1396 <= tmp_ivl_1393 & tmp_ivl_1395;
  LPM_q_ivl_1399 <= tmp_ivl_1401 & tmp_ivl_1396;
  tmp_ivl_1404 <= state_in_s1(303);
  tmp_ivl_1406 <= state_in_s0(303);
  tmp_ivl_1407 <= tmp_ivl_1404 & tmp_ivl_1406;
  LPM_q_ivl_1410 <= tmp_ivl_1412 & tmp_ivl_1407;
  new_AGEMA_signal_2482 <= tmp_ivl_1416(1);
  tmp_ivl_1414 <= tmp_ivl_1416(0);
  tmp_ivl_1416 <= LPM_d0_ivl_1420(0 + 1 downto 0);
  tmp_ivl_1422 <= state_in_s1(302);
  tmp_ivl_1424 <= state_in_s0(302);
  tmp_ivl_1425 <= tmp_ivl_1422 & tmp_ivl_1424;
  LPM_q_ivl_1428 <= tmp_ivl_1430 & tmp_ivl_1425;
  tmp_ivl_1433 <= state_in_s1(238);
  tmp_ivl_1435 <= state_in_s0(238);
  tmp_ivl_1436 <= tmp_ivl_1433 & tmp_ivl_1435;
  LPM_q_ivl_1439 <= tmp_ivl_1441 & tmp_ivl_1436;
  new_AGEMA_signal_2485 <= tmp_ivl_1445(1);
  tmp_ivl_1443 <= tmp_ivl_1445(0);
  tmp_ivl_1445 <= LPM_d0_ivl_1449(0 + 1 downto 0);
  tmp_ivl_1451 <= state_in_s1(301);
  tmp_ivl_1453 <= state_in_s0(301);
  tmp_ivl_1454 <= tmp_ivl_1451 & tmp_ivl_1453;
  LPM_q_ivl_1457 <= tmp_ivl_1459 & tmp_ivl_1454;
  tmp_ivl_1462 <= state_in_s1(237);
  tmp_ivl_1464 <= state_in_s0(237);
  tmp_ivl_1465 <= tmp_ivl_1462 & tmp_ivl_1464;
  LPM_q_ivl_1468 <= tmp_ivl_1470 & tmp_ivl_1465;
  new_AGEMA_signal_2488 <= tmp_ivl_1474(1);
  tmp_ivl_1472 <= tmp_ivl_1474(0);
  tmp_ivl_1474 <= LPM_d0_ivl_1478(0 + 1 downto 0);
  tmp_ivl_1480 <= state_in_s1(236);
  tmp_ivl_1482 <= state_in_s0(236);
  tmp_ivl_1483 <= tmp_ivl_1480 & tmp_ivl_1482;
  LPM_q_ivl_1486 <= tmp_ivl_1488 & tmp_ivl_1483;
  tmp_ivl_1491 <= state_in_s1(300);
  tmp_ivl_1493 <= state_in_s0(300);
  tmp_ivl_1494 <= tmp_ivl_1491 & tmp_ivl_1493;
  LPM_q_ivl_1497 <= tmp_ivl_1499 & tmp_ivl_1494;
  new_AGEMA_signal_2491 <= tmp_ivl_1503(1);
  tmp_ivl_1501 <= tmp_ivl_1503(0);
  tmp_ivl_1503 <= LPM_d0_ivl_1507(0 + 1 downto 0);
  tmp_ivl_1509 <= state_in_s1(313);
  tmp_ivl_1511 <= state_in_s0(313);
  tmp_ivl_1512 <= tmp_ivl_1509 & tmp_ivl_1511;
  LPM_q_ivl_1515 <= tmp_ivl_1517 & tmp_ivl_1512;
  tmp_ivl_1520 <= state_in_s1(249);
  tmp_ivl_1522 <= state_in_s0(249);
  tmp_ivl_1523 <= tmp_ivl_1520 & tmp_ivl_1522;
  LPM_q_ivl_1526 <= tmp_ivl_1528 & tmp_ivl_1523;
  new_AGEMA_signal_2494 <= tmp_ivl_1532(1);
  tmp_ivl_1530 <= tmp_ivl_1532(0);
  tmp_ivl_1532 <= LPM_d0_ivl_1536(0 + 1 downto 0);
  tmp_ivl_1538 <= state_in_s1(235);
  tmp_ivl_1540 <= state_in_s0(235);
  tmp_ivl_1541 <= tmp_ivl_1538 & tmp_ivl_1540;
  LPM_q_ivl_1544 <= tmp_ivl_1546 & tmp_ivl_1541;
  tmp_ivl_1549 <= state_in_s1(299);
  tmp_ivl_1551 <= state_in_s0(299);
  tmp_ivl_1552 <= tmp_ivl_1549 & tmp_ivl_1551;
  LPM_q_ivl_1555 <= tmp_ivl_1557 & tmp_ivl_1552;
  new_AGEMA_signal_2497 <= tmp_ivl_1561(1);
  tmp_ivl_1559 <= tmp_ivl_1561(0);
  tmp_ivl_1561 <= LPM_d0_ivl_1565(0 + 1 downto 0);
  tmp_ivl_1567 <= state_in_s1(298);
  tmp_ivl_1569 <= state_in_s0(298);
  tmp_ivl_1570 <= tmp_ivl_1567 & tmp_ivl_1569;
  LPM_q_ivl_1573 <= tmp_ivl_1575 & tmp_ivl_1570;
  tmp_ivl_1578 <= state_in_s1(234);
  tmp_ivl_1580 <= state_in_s0(234);
  tmp_ivl_1581 <= tmp_ivl_1578 & tmp_ivl_1580;
  LPM_q_ivl_1584 <= tmp_ivl_1586 & tmp_ivl_1581;
  new_AGEMA_signal_2500 <= tmp_ivl_1590(1);
  tmp_ivl_1588 <= tmp_ivl_1590(0);
  tmp_ivl_1590 <= LPM_d0_ivl_1594(0 + 1 downto 0);
  tmp_ivl_1596 <= state_in_s1(233);
  tmp_ivl_1598 <= state_in_s0(233);
  tmp_ivl_1599 <= tmp_ivl_1596 & tmp_ivl_1598;
  LPM_q_ivl_1602 <= tmp_ivl_1604 & tmp_ivl_1599;
  tmp_ivl_1607 <= state_in_s1(297);
  tmp_ivl_1609 <= state_in_s0(297);
  tmp_ivl_1610 <= tmp_ivl_1607 & tmp_ivl_1609;
  LPM_q_ivl_1613 <= tmp_ivl_1615 & tmp_ivl_1610;
  new_AGEMA_signal_2503 <= tmp_ivl_1619(1);
  tmp_ivl_1617 <= tmp_ivl_1619(0);
  tmp_ivl_1619 <= LPM_d0_ivl_1623(0 + 1 downto 0);
  tmp_ivl_1625 <= state_in_s1(232);
  tmp_ivl_1627 <= state_in_s0(232);
  tmp_ivl_1628 <= tmp_ivl_1625 & tmp_ivl_1627;
  LPM_q_ivl_1631 <= tmp_ivl_1633 & tmp_ivl_1628;
  tmp_ivl_1636 <= state_in_s1(296);
  tmp_ivl_1638 <= state_in_s0(296);
  tmp_ivl_1639 <= tmp_ivl_1636 & tmp_ivl_1638;
  LPM_q_ivl_1642 <= tmp_ivl_1644 & tmp_ivl_1639;
  new_AGEMA_signal_2506 <= tmp_ivl_1648(1);
  tmp_ivl_1646 <= tmp_ivl_1648(0);
  tmp_ivl_1648 <= LPM_d0_ivl_1652(0 + 1 downto 0);
  tmp_ivl_1654 <= state_in_s1(311);
  tmp_ivl_1656 <= state_in_s0(311);
  tmp_ivl_1657 <= tmp_ivl_1654 & tmp_ivl_1656;
  LPM_q_ivl_1660 <= tmp_ivl_1662 & tmp_ivl_1657;
  tmp_ivl_1665 <= state_in_s1(247);
  tmp_ivl_1667 <= state_in_s0(247);
  tmp_ivl_1668 <= tmp_ivl_1665 & tmp_ivl_1667;
  LPM_q_ivl_1671 <= tmp_ivl_1673 & tmp_ivl_1668;
  new_AGEMA_signal_2509 <= tmp_ivl_1677(1);
  tmp_ivl_1675 <= tmp_ivl_1677(0);
  tmp_ivl_1677 <= LPM_d0_ivl_1681(0 + 1 downto 0);
  tmp_ivl_1683 <= state_in_s1(246);
  tmp_ivl_1685 <= state_in_s0(246);
  tmp_ivl_1686 <= tmp_ivl_1683 & tmp_ivl_1685;
  LPM_q_ivl_1689 <= tmp_ivl_1691 & tmp_ivl_1686;
  tmp_ivl_1694 <= state_in_s1(310);
  tmp_ivl_1696 <= state_in_s0(310);
  tmp_ivl_1697 <= tmp_ivl_1694 & tmp_ivl_1696;
  LPM_q_ivl_1700 <= tmp_ivl_1702 & tmp_ivl_1697;
  new_AGEMA_signal_2512 <= tmp_ivl_1706(1);
  tmp_ivl_1704 <= tmp_ivl_1706(0);
  tmp_ivl_1706 <= LPM_d0_ivl_1710(0 + 1 downto 0);
  tmp_ivl_1712 <= state_in_s1(245);
  tmp_ivl_1714 <= state_in_s0(245);
  tmp_ivl_1715 <= tmp_ivl_1712 & tmp_ivl_1714;
  LPM_q_ivl_1718 <= tmp_ivl_1720 & tmp_ivl_1715;
  tmp_ivl_1723 <= state_in_s1(309);
  tmp_ivl_1725 <= state_in_s0(309);
  tmp_ivl_1726 <= tmp_ivl_1723 & tmp_ivl_1725;
  LPM_q_ivl_1729 <= tmp_ivl_1731 & tmp_ivl_1726;
  new_AGEMA_signal_2515 <= tmp_ivl_1735(1);
  tmp_ivl_1733 <= tmp_ivl_1735(0);
  tmp_ivl_1735 <= LPM_d0_ivl_1739(0 + 1 downto 0);
  tmp_ivl_1741 <= state_in_s1(244);
  tmp_ivl_1743 <= state_in_s0(244);
  tmp_ivl_1744 <= tmp_ivl_1741 & tmp_ivl_1743;
  LPM_q_ivl_1747 <= tmp_ivl_1749 & tmp_ivl_1744;
  tmp_ivl_1752 <= state_in_s1(308);
  tmp_ivl_1754 <= state_in_s0(308);
  tmp_ivl_1755 <= tmp_ivl_1752 & tmp_ivl_1754;
  LPM_q_ivl_1758 <= tmp_ivl_1760 & tmp_ivl_1755;
  new_AGEMA_signal_2518 <= tmp_ivl_1764(1);
  tmp_ivl_1762 <= tmp_ivl_1764(0);
  tmp_ivl_1764 <= LPM_d0_ivl_1768(0 + 1 downto 0);
  tmp_ivl_1770 <= state_in_s1(307);
  tmp_ivl_1772 <= state_in_s0(307);
  tmp_ivl_1773 <= tmp_ivl_1770 & tmp_ivl_1772;
  LPM_q_ivl_1776 <= tmp_ivl_1778 & tmp_ivl_1773;
  tmp_ivl_1781 <= state_in_s1(243);
  tmp_ivl_1783 <= state_in_s0(243);
  tmp_ivl_1784 <= tmp_ivl_1781 & tmp_ivl_1783;
  LPM_q_ivl_1787 <= tmp_ivl_1789 & tmp_ivl_1784;
  new_AGEMA_signal_2521 <= tmp_ivl_1793(1);
  tmp_ivl_1791 <= tmp_ivl_1793(0);
  tmp_ivl_1793 <= LPM_d0_ivl_1797(0 + 1 downto 0);
  tmp_ivl_1799 <= state_in_s1(242);
  tmp_ivl_1801 <= state_in_s0(242);
  tmp_ivl_1802 <= tmp_ivl_1799 & tmp_ivl_1801;
  LPM_q_ivl_1805 <= tmp_ivl_1807 & tmp_ivl_1802;
  tmp_ivl_1810 <= state_in_s1(306);
  tmp_ivl_1812 <= state_in_s0(306);
  tmp_ivl_1813 <= tmp_ivl_1810 & tmp_ivl_1812;
  LPM_q_ivl_1816 <= tmp_ivl_1818 & tmp_ivl_1813;
  new_AGEMA_signal_2524 <= tmp_ivl_1822(1);
  tmp_ivl_1820 <= tmp_ivl_1822(0);
  tmp_ivl_1822 <= LPM_d0_ivl_1826(0 + 1 downto 0);
  tmp_ivl_1828 <= state_in_s1(248);
  tmp_ivl_1830 <= state_in_s0(248);
  tmp_ivl_1831 <= tmp_ivl_1828 & tmp_ivl_1830;
  LPM_q_ivl_1834 <= tmp_ivl_1836 & tmp_ivl_1831;
  tmp_ivl_1839 <= state_in_s1(312);
  tmp_ivl_1841 <= state_in_s0(312);
  tmp_ivl_1842 <= tmp_ivl_1839 & tmp_ivl_1841;
  LPM_q_ivl_1845 <= tmp_ivl_1847 & tmp_ivl_1842;
  new_AGEMA_signal_2527 <= tmp_ivl_1851(1);
  tmp_ivl_1849 <= tmp_ivl_1851(0);
  tmp_ivl_1851 <= LPM_d0_ivl_1855(0 + 1 downto 0);
  tmp_ivl_1857 <= state_in_s1(49);
  tmp_ivl_1859 <= state_in_s0(49);
  tmp_ivl_1860 <= tmp_ivl_1857 & tmp_ivl_1859;
  LPM_q_ivl_1863 <= tmp_ivl_1865 & tmp_ivl_1860;
  tmp_ivl_1868 <= state_in_s1(305);
  tmp_ivl_1870 <= state_in_s0(305);
  tmp_ivl_1871 <= tmp_ivl_1868 & tmp_ivl_1870;
  LPM_q_ivl_1874 <= tmp_ivl_1876 & tmp_ivl_1871;
  new_AGEMA_signal_2529 <= tmp_ivl_1880(1);
  tmp_ivl_1878 <= tmp_ivl_1880(0);
  tmp_ivl_1880 <= LPM_d0_ivl_1884(0 + 1 downto 0);
  tmp_ivl_1886 <= state_in_s1(48);
  tmp_ivl_1888 <= state_in_s0(48);
  tmp_ivl_1889 <= tmp_ivl_1886 & tmp_ivl_1888;
  LPM_q_ivl_1892 <= tmp_ivl_1894 & tmp_ivl_1889;
  tmp_ivl_1897 <= state_in_s1(304);
  tmp_ivl_1899 <= state_in_s0(304);
  tmp_ivl_1900 <= tmp_ivl_1897 & tmp_ivl_1899;
  LPM_q_ivl_1903 <= tmp_ivl_1905 & tmp_ivl_1900;
  new_AGEMA_signal_2531 <= tmp_ivl_1909(1);
  tmp_ivl_1907 <= tmp_ivl_1909(0);
  tmp_ivl_1909 <= LPM_d0_ivl_1913(0 + 1 downto 0);
  tmp_ivl_1915 <= state_in_s1(63);
  tmp_ivl_1917 <= state_in_s0(63);
  tmp_ivl_1918 <= tmp_ivl_1915 & tmp_ivl_1917;
  LPM_q_ivl_1921 <= tmp_ivl_1923 & tmp_ivl_1918;
  tmp_ivl_1926 <= state_in_s1(319);
  tmp_ivl_1928 <= state_in_s0(319);
  tmp_ivl_1929 <= tmp_ivl_1926 & tmp_ivl_1928;
  LPM_q_ivl_1932 <= tmp_ivl_1934 & tmp_ivl_1929;
  new_AGEMA_signal_2533 <= tmp_ivl_1938(1);
  tmp_ivl_1936 <= tmp_ivl_1938(0);
  tmp_ivl_1938 <= LPM_d0_ivl_1942(0 + 1 downto 0);
  tmp_ivl_1944 <= state_in_s1(62);
  tmp_ivl_1946 <= state_in_s0(62);
  tmp_ivl_1947 <= tmp_ivl_1944 & tmp_ivl_1946;
  LPM_q_ivl_1950 <= tmp_ivl_1952 & tmp_ivl_1947;
  tmp_ivl_1955 <= state_in_s1(318);
  tmp_ivl_1957 <= state_in_s0(318);
  tmp_ivl_1958 <= tmp_ivl_1955 & tmp_ivl_1957;
  LPM_q_ivl_1961 <= tmp_ivl_1963 & tmp_ivl_1958;
  new_AGEMA_signal_2535 <= tmp_ivl_1967(1);
  tmp_ivl_1965 <= tmp_ivl_1967(0);
  tmp_ivl_1967 <= LPM_d0_ivl_1971(0 + 1 downto 0);
  tmp_ivl_1973 <= state_in_s1(7);
  tmp_ivl_1975 <= state_in_s0(7);
  tmp_ivl_1976 <= tmp_ivl_1973 & tmp_ivl_1975;
  LPM_q_ivl_1979 <= tmp_ivl_1981 & tmp_ivl_1976;
  tmp_ivl_1984 <= state_in_s1(263);
  tmp_ivl_1986 <= state_in_s0(263);
  tmp_ivl_1987 <= tmp_ivl_1984 & tmp_ivl_1986;
  LPM_q_ivl_1990 <= tmp_ivl_1992 & tmp_ivl_1987;
  new_AGEMA_signal_2537 <= tmp_ivl_1996(1);
  tmp_ivl_1994 <= tmp_ivl_1996(0);
  tmp_ivl_1996 <= LPM_d0_ivl_2000(0 + 1 downto 0);
  tmp_ivl_2002 <= state_in_s1(6);
  tmp_ivl_2004 <= state_in_s0(6);
  tmp_ivl_2005 <= tmp_ivl_2002 & tmp_ivl_2004;
  LPM_q_ivl_2008 <= tmp_ivl_2010 & tmp_ivl_2005;
  tmp_ivl_2013 <= state_in_s1(262);
  tmp_ivl_2015 <= state_in_s0(262);
  tmp_ivl_2016 <= tmp_ivl_2013 & tmp_ivl_2015;
  LPM_q_ivl_2019 <= tmp_ivl_2021 & tmp_ivl_2016;
  new_AGEMA_signal_2539 <= tmp_ivl_2025(1);
  tmp_ivl_2023 <= tmp_ivl_2025(0);
  tmp_ivl_2025 <= LPM_d0_ivl_2029(0 + 1 downto 0);
  tmp_ivl_2031 <= state_in_s1(5);
  tmp_ivl_2033 <= state_in_s0(5);
  tmp_ivl_2034 <= tmp_ivl_2031 & tmp_ivl_2033;
  LPM_q_ivl_2037 <= tmp_ivl_2039 & tmp_ivl_2034;
  tmp_ivl_2042 <= state_in_s1(261);
  tmp_ivl_2044 <= state_in_s0(261);
  tmp_ivl_2045 <= tmp_ivl_2042 & tmp_ivl_2044;
  LPM_q_ivl_2048 <= tmp_ivl_2050 & tmp_ivl_2045;
  new_AGEMA_signal_2541 <= tmp_ivl_2054(1);
  tmp_ivl_2052 <= tmp_ivl_2054(0);
  tmp_ivl_2054 <= LPM_d0_ivl_2058(0 + 1 downto 0);
  tmp_ivl_2060 <= state_in_s1(4);
  tmp_ivl_2062 <= state_in_s0(4);
  tmp_ivl_2063 <= tmp_ivl_2060 & tmp_ivl_2062;
  LPM_q_ivl_2066 <= tmp_ivl_2068 & tmp_ivl_2063;
  tmp_ivl_2071 <= state_in_s1(260);
  tmp_ivl_2073 <= state_in_s0(260);
  tmp_ivl_2074 <= tmp_ivl_2071 & tmp_ivl_2073;
  LPM_q_ivl_2077 <= tmp_ivl_2079 & tmp_ivl_2074;
  new_AGEMA_signal_2543 <= tmp_ivl_2083(1);
  tmp_ivl_2081 <= tmp_ivl_2083(0);
  tmp_ivl_2083 <= LPM_d0_ivl_2087(0 + 1 downto 0);
  tmp_ivl_2089 <= state_in_s1(61);
  tmp_ivl_2091 <= state_in_s0(61);
  tmp_ivl_2092 <= tmp_ivl_2089 & tmp_ivl_2091;
  LPM_q_ivl_2095 <= tmp_ivl_2097 & tmp_ivl_2092;
  tmp_ivl_2100 <= state_in_s1(317);
  tmp_ivl_2102 <= state_in_s0(317);
  tmp_ivl_2103 <= tmp_ivl_2100 & tmp_ivl_2102;
  LPM_q_ivl_2106 <= tmp_ivl_2108 & tmp_ivl_2103;
  new_AGEMA_signal_2545 <= tmp_ivl_2112(1);
  tmp_ivl_2110 <= tmp_ivl_2112(0);
  tmp_ivl_2112 <= LPM_d0_ivl_2116(0 + 1 downto 0);
  tmp_ivl_2118 <= state_in_s1(259);
  tmp_ivl_2120 <= state_in_s0(259);
  tmp_ivl_2121 <= tmp_ivl_2118 & tmp_ivl_2120;
  LPM_q_ivl_2124 <= tmp_ivl_2126 & tmp_ivl_2121;
  tmp_ivl_2129 <= state_in_s1(3);
  tmp_ivl_2131 <= state_in_s0(3);
  tmp_ivl_2132 <= tmp_ivl_2129 & tmp_ivl_2131;
  LPM_q_ivl_2135 <= tmp_ivl_2137 & tmp_ivl_2132;
  new_AGEMA_signal_2547 <= tmp_ivl_2141(1);
  tmp_ivl_2139 <= tmp_ivl_2141(0);
  tmp_ivl_2141 <= LPM_d0_ivl_2145(0 + 1 downto 0);
  tmp_ivl_2147 <= state_in_s1(258);
  tmp_ivl_2149 <= state_in_s0(258);
  tmp_ivl_2150 <= tmp_ivl_2147 & tmp_ivl_2149;
  LPM_q_ivl_2153 <= tmp_ivl_2155 & tmp_ivl_2150;
  tmp_ivl_2158 <= state_in_s1(2);
  tmp_ivl_2160 <= state_in_s0(2);
  tmp_ivl_2161 <= tmp_ivl_2158 & tmp_ivl_2160;
  LPM_q_ivl_2164 <= tmp_ivl_2166 & tmp_ivl_2161;
  new_AGEMA_signal_2549 <= tmp_ivl_2170(1);
  tmp_ivl_2168 <= tmp_ivl_2170(0);
  tmp_ivl_2170 <= LPM_d0_ivl_2174(0 + 1 downto 0);
  tmp_ivl_2176 <= state_in_s1(257);
  tmp_ivl_2178 <= state_in_s0(257);
  tmp_ivl_2179 <= tmp_ivl_2176 & tmp_ivl_2178;
  LPM_q_ivl_2182 <= tmp_ivl_2184 & tmp_ivl_2179;
  tmp_ivl_2187 <= state_in_s1(1);
  tmp_ivl_2189 <= state_in_s0(1);
  tmp_ivl_2190 <= tmp_ivl_2187 & tmp_ivl_2189;
  LPM_q_ivl_2193 <= tmp_ivl_2195 & tmp_ivl_2190;
  new_AGEMA_signal_2551 <= tmp_ivl_2199(1);
  tmp_ivl_2197 <= tmp_ivl_2199(0);
  tmp_ivl_2199 <= LPM_d0_ivl_2203(0 + 1 downto 0);
  tmp_ivl_2205 <= state_in_s1(0);
  tmp_ivl_2207 <= state_in_s0(0);
  tmp_ivl_2208 <= tmp_ivl_2205 & tmp_ivl_2207;
  LPM_q_ivl_2211 <= tmp_ivl_2213 & tmp_ivl_2208;
  tmp_ivl_2216 <= state_in_s1(256);
  tmp_ivl_2218 <= state_in_s0(256);
  tmp_ivl_2219 <= tmp_ivl_2216 & tmp_ivl_2218;
  LPM_q_ivl_2222 <= tmp_ivl_2224 & tmp_ivl_2219;
  new_AGEMA_signal_2553 <= tmp_ivl_2228(1);
  tmp_ivl_2226 <= tmp_ivl_2228(0);
  tmp_ivl_2228 <= LPM_d0_ivl_2232(0 + 1 downto 0);
  tmp_ivl_2234 <= state_in_s1(15);
  tmp_ivl_2236 <= state_in_s0(15);
  tmp_ivl_2237 <= tmp_ivl_2234 & tmp_ivl_2236;
  LPM_q_ivl_2240 <= tmp_ivl_2242 & tmp_ivl_2237;
  tmp_ivl_2245 <= state_in_s1(271);
  tmp_ivl_2247 <= state_in_s0(271);
  tmp_ivl_2248 <= tmp_ivl_2245 & tmp_ivl_2247;
  LPM_q_ivl_2251 <= tmp_ivl_2253 & tmp_ivl_2248;
  new_AGEMA_signal_2555 <= tmp_ivl_2257(1);
  tmp_ivl_2255 <= tmp_ivl_2257(0);
  tmp_ivl_2257 <= LPM_d0_ivl_2261(0 + 1 downto 0);
  tmp_ivl_2263 <= state_in_s1(14);
  tmp_ivl_2265 <= state_in_s0(14);
  tmp_ivl_2266 <= tmp_ivl_2263 & tmp_ivl_2265;
  LPM_q_ivl_2269 <= tmp_ivl_2271 & tmp_ivl_2266;
  tmp_ivl_2274 <= state_in_s1(270);
  tmp_ivl_2276 <= state_in_s0(270);
  tmp_ivl_2277 <= tmp_ivl_2274 & tmp_ivl_2276;
  LPM_q_ivl_2280 <= tmp_ivl_2282 & tmp_ivl_2277;
  new_AGEMA_signal_2557 <= tmp_ivl_2286(1);
  tmp_ivl_2284 <= tmp_ivl_2286(0);
  tmp_ivl_2286 <= LPM_d0_ivl_2290(0 + 1 downto 0);
  tmp_ivl_2292 <= state_in_s1(13);
  tmp_ivl_2294 <= state_in_s0(13);
  tmp_ivl_2295 <= tmp_ivl_2292 & tmp_ivl_2294;
  LPM_q_ivl_2298 <= tmp_ivl_2300 & tmp_ivl_2295;
  tmp_ivl_2303 <= state_in_s1(269);
  tmp_ivl_2305 <= state_in_s0(269);
  tmp_ivl_2306 <= tmp_ivl_2303 & tmp_ivl_2305;
  LPM_q_ivl_2309 <= tmp_ivl_2311 & tmp_ivl_2306;
  new_AGEMA_signal_2559 <= tmp_ivl_2315(1);
  tmp_ivl_2313 <= tmp_ivl_2315(0);
  tmp_ivl_2315 <= LPM_d0_ivl_2319(0 + 1 downto 0);
  tmp_ivl_2321 <= state_in_s1(268);
  tmp_ivl_2323 <= state_in_s0(268);
  tmp_ivl_2324 <= tmp_ivl_2321 & tmp_ivl_2323;
  LPM_q_ivl_2327 <= tmp_ivl_2329 & tmp_ivl_2324;
  tmp_ivl_2332 <= state_in_s1(12);
  tmp_ivl_2334 <= state_in_s0(12);
  tmp_ivl_2335 <= tmp_ivl_2332 & tmp_ivl_2334;
  LPM_q_ivl_2338 <= tmp_ivl_2340 & tmp_ivl_2335;
  new_AGEMA_signal_2561 <= tmp_ivl_2344(1);
  tmp_ivl_2342 <= tmp_ivl_2344(0);
  tmp_ivl_2344 <= LPM_d0_ivl_2348(0 + 1 downto 0);
  tmp_ivl_2350 <= state_in_s1(267);
  tmp_ivl_2352 <= state_in_s0(267);
  tmp_ivl_2353 <= tmp_ivl_2350 & tmp_ivl_2352;
  LPM_q_ivl_2356 <= tmp_ivl_2358 & tmp_ivl_2353;
  tmp_ivl_2361 <= state_in_s1(11);
  tmp_ivl_2363 <= state_in_s0(11);
  tmp_ivl_2364 <= tmp_ivl_2361 & tmp_ivl_2363;
  LPM_q_ivl_2367 <= tmp_ivl_2369 & tmp_ivl_2364;
  new_AGEMA_signal_2563 <= tmp_ivl_2373(1);
  tmp_ivl_2371 <= tmp_ivl_2373(0);
  tmp_ivl_2373 <= LPM_d0_ivl_2377(0 + 1 downto 0);
  tmp_ivl_2379 <= state_in_s1(10);
  tmp_ivl_2381 <= state_in_s0(10);
  tmp_ivl_2382 <= tmp_ivl_2379 & tmp_ivl_2381;
  LPM_q_ivl_2385 <= tmp_ivl_2387 & tmp_ivl_2382;
  tmp_ivl_2390 <= state_in_s1(266);
  tmp_ivl_2392 <= state_in_s0(266);
  tmp_ivl_2393 <= tmp_ivl_2390 & tmp_ivl_2392;
  LPM_q_ivl_2396 <= tmp_ivl_2398 & tmp_ivl_2393;
  new_AGEMA_signal_2565 <= tmp_ivl_2402(1);
  tmp_ivl_2400 <= tmp_ivl_2402(0);
  tmp_ivl_2402 <= LPM_d0_ivl_2406(0 + 1 downto 0);
  tmp_ivl_2408 <= state_in_s1(60);
  tmp_ivl_2410 <= state_in_s0(60);
  tmp_ivl_2411 <= tmp_ivl_2408 & tmp_ivl_2410;
  LPM_q_ivl_2414 <= tmp_ivl_2416 & tmp_ivl_2411;
  tmp_ivl_2419 <= state_in_s1(316);
  tmp_ivl_2421 <= state_in_s0(316);
  tmp_ivl_2422 <= tmp_ivl_2419 & tmp_ivl_2421;
  LPM_q_ivl_2425 <= tmp_ivl_2427 & tmp_ivl_2422;
  new_AGEMA_signal_2567 <= tmp_ivl_2431(1);
  tmp_ivl_2429 <= tmp_ivl_2431(0);
  tmp_ivl_2431 <= LPM_d0_ivl_2435(0 + 1 downto 0);
  tmp_ivl_2437 <= state_in_s1(9);
  tmp_ivl_2439 <= state_in_s0(9);
  tmp_ivl_2440 <= tmp_ivl_2437 & tmp_ivl_2439;
  LPM_q_ivl_2443 <= tmp_ivl_2445 & tmp_ivl_2440;
  tmp_ivl_2448 <= state_in_s1(265);
  tmp_ivl_2450 <= state_in_s0(265);
  tmp_ivl_2451 <= tmp_ivl_2448 & tmp_ivl_2450;
  LPM_q_ivl_2454 <= tmp_ivl_2456 & tmp_ivl_2451;
  new_AGEMA_signal_2569 <= tmp_ivl_2460(1);
  tmp_ivl_2458 <= tmp_ivl_2460(0);
  tmp_ivl_2460 <= LPM_d0_ivl_2464(0 + 1 downto 0);
  tmp_ivl_2466 <= state_in_s1(264);
  tmp_ivl_2468 <= state_in_s0(264);
  tmp_ivl_2469 <= tmp_ivl_2466 & tmp_ivl_2468;
  LPM_q_ivl_2472 <= tmp_ivl_2474 & tmp_ivl_2469;
  tmp_ivl_2477 <= state_in_s1(8);
  tmp_ivl_2479 <= state_in_s0(8);
  tmp_ivl_2480 <= tmp_ivl_2477 & tmp_ivl_2479;
  LPM_q_ivl_2483 <= tmp_ivl_2485 & tmp_ivl_2480;
  new_AGEMA_signal_2571 <= tmp_ivl_2489(1);
  tmp_ivl_2487 <= tmp_ivl_2489(0);
  tmp_ivl_2489 <= LPM_d0_ivl_2493(0 + 1 downto 0);
  tmp_ivl_2495 <= state_in_s1(279);
  tmp_ivl_2497 <= state_in_s0(279);
  tmp_ivl_2498 <= tmp_ivl_2495 & tmp_ivl_2497;
  LPM_q_ivl_2501 <= tmp_ivl_2503 & tmp_ivl_2498;
  tmp_ivl_2506 <= state_in_s1(23);
  tmp_ivl_2508 <= state_in_s0(23);
  tmp_ivl_2509 <= tmp_ivl_2506 & tmp_ivl_2508;
  LPM_q_ivl_2512 <= tmp_ivl_2514 & tmp_ivl_2509;
  new_AGEMA_signal_2573 <= tmp_ivl_2518(1);
  tmp_ivl_2516 <= tmp_ivl_2518(0);
  tmp_ivl_2518 <= LPM_d0_ivl_2522(0 + 1 downto 0);
  tmp_ivl_2524 <= state_in_s1(22);
  tmp_ivl_2526 <= state_in_s0(22);
  tmp_ivl_2527 <= tmp_ivl_2524 & tmp_ivl_2526;
  LPM_q_ivl_2530 <= tmp_ivl_2532 & tmp_ivl_2527;
  tmp_ivl_2535 <= state_in_s1(278);
  tmp_ivl_2537 <= state_in_s0(278);
  tmp_ivl_2538 <= tmp_ivl_2535 & tmp_ivl_2537;
  LPM_q_ivl_2541 <= tmp_ivl_2543 & tmp_ivl_2538;
  new_AGEMA_signal_2575 <= tmp_ivl_2547(1);
  tmp_ivl_2545 <= tmp_ivl_2547(0);
  tmp_ivl_2547 <= LPM_d0_ivl_2551(0 + 1 downto 0);
  tmp_ivl_2553 <= state_in_s1(277);
  tmp_ivl_2555 <= state_in_s0(277);
  tmp_ivl_2556 <= tmp_ivl_2553 & tmp_ivl_2555;
  LPM_q_ivl_2559 <= tmp_ivl_2561 & tmp_ivl_2556;
  tmp_ivl_2564 <= state_in_s1(21);
  tmp_ivl_2566 <= state_in_s0(21);
  tmp_ivl_2567 <= tmp_ivl_2564 & tmp_ivl_2566;
  LPM_q_ivl_2570 <= tmp_ivl_2572 & tmp_ivl_2567;
  new_AGEMA_signal_2577 <= tmp_ivl_2576(1);
  tmp_ivl_2574 <= tmp_ivl_2576(0);
  tmp_ivl_2576 <= LPM_d0_ivl_2580(0 + 1 downto 0);
  tmp_ivl_2582 <= state_in_s1(276);
  tmp_ivl_2584 <= state_in_s0(276);
  tmp_ivl_2585 <= tmp_ivl_2582 & tmp_ivl_2584;
  LPM_q_ivl_2588 <= tmp_ivl_2590 & tmp_ivl_2585;
  tmp_ivl_2593 <= state_in_s1(20);
  tmp_ivl_2595 <= state_in_s0(20);
  tmp_ivl_2596 <= tmp_ivl_2593 & tmp_ivl_2595;
  LPM_q_ivl_2599 <= tmp_ivl_2601 & tmp_ivl_2596;
  new_AGEMA_signal_2579 <= tmp_ivl_2605(1);
  tmp_ivl_2603 <= tmp_ivl_2605(0);
  tmp_ivl_2605 <= LPM_d0_ivl_2609(0 + 1 downto 0);
  tmp_ivl_2611 <= state_in_s1(19);
  tmp_ivl_2613 <= state_in_s0(19);
  tmp_ivl_2614 <= tmp_ivl_2611 & tmp_ivl_2613;
  LPM_q_ivl_2617 <= tmp_ivl_2619 & tmp_ivl_2614;
  tmp_ivl_2622 <= state_in_s1(275);
  tmp_ivl_2624 <= state_in_s0(275);
  tmp_ivl_2625 <= tmp_ivl_2622 & tmp_ivl_2624;
  LPM_q_ivl_2628 <= tmp_ivl_2630 & tmp_ivl_2625;
  new_AGEMA_signal_2581 <= tmp_ivl_2634(1);
  tmp_ivl_2632 <= tmp_ivl_2634(0);
  tmp_ivl_2634 <= LPM_d0_ivl_2638(0 + 1 downto 0);
  tmp_ivl_2640 <= state_in_s1(18);
  tmp_ivl_2642 <= state_in_s0(18);
  tmp_ivl_2643 <= tmp_ivl_2640 & tmp_ivl_2642;
  LPM_q_ivl_2646 <= tmp_ivl_2648 & tmp_ivl_2643;
  tmp_ivl_2651 <= state_in_s1(274);
  tmp_ivl_2653 <= state_in_s0(274);
  tmp_ivl_2654 <= tmp_ivl_2651 & tmp_ivl_2653;
  LPM_q_ivl_2657 <= tmp_ivl_2659 & tmp_ivl_2654;
  new_AGEMA_signal_2583 <= tmp_ivl_2663(1);
  tmp_ivl_2661 <= tmp_ivl_2663(0);
  tmp_ivl_2663 <= LPM_d0_ivl_2667(0 + 1 downto 0);
  tmp_ivl_2669 <= state_in_s1(273);
  tmp_ivl_2671 <= state_in_s0(273);
  tmp_ivl_2672 <= tmp_ivl_2669 & tmp_ivl_2671;
  LPM_q_ivl_2675 <= tmp_ivl_2677 & tmp_ivl_2672;
  tmp_ivl_2680 <= state_in_s1(17);
  tmp_ivl_2682 <= state_in_s0(17);
  tmp_ivl_2683 <= tmp_ivl_2680 & tmp_ivl_2682;
  LPM_q_ivl_2686 <= tmp_ivl_2688 & tmp_ivl_2683;
  new_AGEMA_signal_2585 <= tmp_ivl_2692(1);
  tmp_ivl_2690 <= tmp_ivl_2692(0);
  tmp_ivl_2692 <= LPM_d0_ivl_2696(0 + 1 downto 0);
  tmp_ivl_2698 <= state_in_s1(16);
  tmp_ivl_2700 <= state_in_s0(16);
  tmp_ivl_2701 <= tmp_ivl_2698 & tmp_ivl_2700;
  LPM_q_ivl_2704 <= tmp_ivl_2706 & tmp_ivl_2701;
  tmp_ivl_2709 <= state_in_s1(272);
  tmp_ivl_2711 <= state_in_s0(272);
  tmp_ivl_2712 <= tmp_ivl_2709 & tmp_ivl_2711;
  LPM_q_ivl_2715 <= tmp_ivl_2717 & tmp_ivl_2712;
  new_AGEMA_signal_2587 <= tmp_ivl_2721(1);
  tmp_ivl_2719 <= tmp_ivl_2721(0);
  tmp_ivl_2721 <= LPM_d0_ivl_2725(0 + 1 downto 0);
  tmp_ivl_2727 <= state_in_s1(59);
  tmp_ivl_2729 <= state_in_s0(59);
  tmp_ivl_2730 <= tmp_ivl_2727 & tmp_ivl_2729;
  LPM_q_ivl_2733 <= tmp_ivl_2735 & tmp_ivl_2730;
  tmp_ivl_2738 <= state_in_s1(315);
  tmp_ivl_2740 <= state_in_s0(315);
  tmp_ivl_2741 <= tmp_ivl_2738 & tmp_ivl_2740;
  LPM_q_ivl_2744 <= tmp_ivl_2746 & tmp_ivl_2741;
  new_AGEMA_signal_2589 <= tmp_ivl_2750(1);
  tmp_ivl_2748 <= tmp_ivl_2750(0);
  tmp_ivl_2750 <= LPM_d0_ivl_2754(0 + 1 downto 0);
  tmp_ivl_2756 <= state_in_s1(31);
  tmp_ivl_2758 <= state_in_s0(31);
  tmp_ivl_2759 <= tmp_ivl_2756 & tmp_ivl_2758;
  LPM_q_ivl_2762 <= tmp_ivl_2764 & tmp_ivl_2759;
  tmp_ivl_2767 <= state_in_s1(287);
  tmp_ivl_2769 <= state_in_s0(287);
  tmp_ivl_2770 <= tmp_ivl_2767 & tmp_ivl_2769;
  LPM_q_ivl_2773 <= tmp_ivl_2775 & tmp_ivl_2770;
  new_AGEMA_signal_2591 <= tmp_ivl_2779(1);
  tmp_ivl_2777 <= tmp_ivl_2779(0);
  tmp_ivl_2779 <= LPM_d0_ivl_2783(0 + 1 downto 0);
  tmp_ivl_2785 <= state_in_s1(30);
  tmp_ivl_2787 <= state_in_s0(30);
  tmp_ivl_2788 <= tmp_ivl_2785 & tmp_ivl_2787;
  LPM_q_ivl_2791 <= tmp_ivl_2793 & tmp_ivl_2788;
  tmp_ivl_2796 <= state_in_s1(286);
  tmp_ivl_2798 <= state_in_s0(286);
  tmp_ivl_2799 <= tmp_ivl_2796 & tmp_ivl_2798;
  LPM_q_ivl_2802 <= tmp_ivl_2804 & tmp_ivl_2799;
  new_AGEMA_signal_2593 <= tmp_ivl_2808(1);
  tmp_ivl_2806 <= tmp_ivl_2808(0);
  tmp_ivl_2808 <= LPM_d0_ivl_2812(0 + 1 downto 0);
  tmp_ivl_2814 <= state_in_s1(29);
  tmp_ivl_2816 <= state_in_s0(29);
  tmp_ivl_2817 <= tmp_ivl_2814 & tmp_ivl_2816;
  LPM_q_ivl_2820 <= tmp_ivl_2822 & tmp_ivl_2817;
  tmp_ivl_2825 <= state_in_s1(285);
  tmp_ivl_2827 <= state_in_s0(285);
  tmp_ivl_2828 <= tmp_ivl_2825 & tmp_ivl_2827;
  LPM_q_ivl_2831 <= tmp_ivl_2833 & tmp_ivl_2828;
  new_AGEMA_signal_2595 <= tmp_ivl_2837(1);
  tmp_ivl_2835 <= tmp_ivl_2837(0);
  tmp_ivl_2837 <= LPM_d0_ivl_2841(0 + 1 downto 0);
  tmp_ivl_2843 <= state_in_s1(28);
  tmp_ivl_2845 <= state_in_s0(28);
  tmp_ivl_2846 <= tmp_ivl_2843 & tmp_ivl_2845;
  LPM_q_ivl_2849 <= tmp_ivl_2851 & tmp_ivl_2846;
  tmp_ivl_2854 <= state_in_s1(284);
  tmp_ivl_2856 <= state_in_s0(284);
  tmp_ivl_2857 <= tmp_ivl_2854 & tmp_ivl_2856;
  LPM_q_ivl_2860 <= tmp_ivl_2862 & tmp_ivl_2857;
  new_AGEMA_signal_2597 <= tmp_ivl_2866(1);
  tmp_ivl_2864 <= tmp_ivl_2866(0);
  tmp_ivl_2866 <= LPM_d0_ivl_2870(0 + 1 downto 0);
  tmp_ivl_2872 <= state_in_s1(27);
  tmp_ivl_2874 <= state_in_s0(27);
  tmp_ivl_2875 <= tmp_ivl_2872 & tmp_ivl_2874;
  LPM_q_ivl_2878 <= tmp_ivl_2880 & tmp_ivl_2875;
  tmp_ivl_2883 <= state_in_s1(283);
  tmp_ivl_2885 <= state_in_s0(283);
  tmp_ivl_2886 <= tmp_ivl_2883 & tmp_ivl_2885;
  LPM_q_ivl_2889 <= tmp_ivl_2891 & tmp_ivl_2886;
  new_AGEMA_signal_2599 <= tmp_ivl_2895(1);
  tmp_ivl_2893 <= tmp_ivl_2895(0);
  tmp_ivl_2895 <= LPM_d0_ivl_2899(0 + 1 downto 0);
  tmp_ivl_2901 <= state_in_s1(26);
  tmp_ivl_2903 <= state_in_s0(26);
  tmp_ivl_2904 <= tmp_ivl_2901 & tmp_ivl_2903;
  LPM_q_ivl_2907 <= tmp_ivl_2909 & tmp_ivl_2904;
  tmp_ivl_2912 <= state_in_s1(282);
  tmp_ivl_2914 <= state_in_s0(282);
  tmp_ivl_2915 <= tmp_ivl_2912 & tmp_ivl_2914;
  LPM_q_ivl_2918 <= tmp_ivl_2920 & tmp_ivl_2915;
  new_AGEMA_signal_2601 <= tmp_ivl_2924(1);
  tmp_ivl_2922 <= tmp_ivl_2924(0);
  tmp_ivl_2924 <= LPM_d0_ivl_2928(0 + 1 downto 0);
  tmp_ivl_2930 <= state_in_s1(25);
  tmp_ivl_2932 <= state_in_s0(25);
  tmp_ivl_2933 <= tmp_ivl_2930 & tmp_ivl_2932;
  LPM_q_ivl_2936 <= tmp_ivl_2938 & tmp_ivl_2933;
  tmp_ivl_2941 <= state_in_s1(281);
  tmp_ivl_2943 <= state_in_s0(281);
  tmp_ivl_2944 <= tmp_ivl_2941 & tmp_ivl_2943;
  LPM_q_ivl_2947 <= tmp_ivl_2949 & tmp_ivl_2944;
  new_AGEMA_signal_2603 <= tmp_ivl_2953(1);
  tmp_ivl_2951 <= tmp_ivl_2953(0);
  tmp_ivl_2953 <= LPM_d0_ivl_2957(0 + 1 downto 0);
  tmp_ivl_2959 <= state_in_s1(24);
  tmp_ivl_2961 <= state_in_s0(24);
  tmp_ivl_2962 <= tmp_ivl_2959 & tmp_ivl_2961;
  LPM_q_ivl_2965 <= tmp_ivl_2967 & tmp_ivl_2962;
  tmp_ivl_2970 <= state_in_s1(280);
  tmp_ivl_2972 <= state_in_s0(280);
  tmp_ivl_2973 <= tmp_ivl_2970 & tmp_ivl_2972;
  LPM_q_ivl_2976 <= tmp_ivl_2978 & tmp_ivl_2973;
  new_AGEMA_signal_2605 <= tmp_ivl_2982(1);
  tmp_ivl_2980 <= tmp_ivl_2982(0);
  tmp_ivl_2982 <= LPM_d0_ivl_2986(0 + 1 downto 0);
  tmp_ivl_2988 <= state_in_s1(39);
  tmp_ivl_2990 <= state_in_s0(39);
  tmp_ivl_2991 <= tmp_ivl_2988 & tmp_ivl_2990;
  LPM_q_ivl_2994 <= tmp_ivl_2996 & tmp_ivl_2991;
  tmp_ivl_2999 <= state_in_s1(295);
  tmp_ivl_3001 <= state_in_s0(295);
  tmp_ivl_3002 <= tmp_ivl_2999 & tmp_ivl_3001;
  LPM_q_ivl_3005 <= tmp_ivl_3007 & tmp_ivl_3002;
  new_AGEMA_signal_2607 <= tmp_ivl_3011(1);
  tmp_ivl_3009 <= tmp_ivl_3011(0);
  tmp_ivl_3011 <= LPM_d0_ivl_3015(0 + 1 downto 0);
  tmp_ivl_3017 <= state_in_s1(38);
  tmp_ivl_3019 <= state_in_s0(38);
  tmp_ivl_3020 <= tmp_ivl_3017 & tmp_ivl_3019;
  LPM_q_ivl_3023 <= tmp_ivl_3025 & tmp_ivl_3020;
  tmp_ivl_3028 <= state_in_s1(294);
  tmp_ivl_3030 <= state_in_s0(294);
  tmp_ivl_3031 <= tmp_ivl_3028 & tmp_ivl_3030;
  LPM_q_ivl_3034 <= tmp_ivl_3036 & tmp_ivl_3031;
  new_AGEMA_signal_2609 <= tmp_ivl_3040(1);
  tmp_ivl_3038 <= tmp_ivl_3040(0);
  tmp_ivl_3040 <= LPM_d0_ivl_3044(0 + 1 downto 0);
  tmp_ivl_3046 <= state_in_s1(58);
  tmp_ivl_3048 <= state_in_s0(58);
  tmp_ivl_3049 <= tmp_ivl_3046 & tmp_ivl_3048;
  LPM_q_ivl_3052 <= tmp_ivl_3054 & tmp_ivl_3049;
  tmp_ivl_3057 <= state_in_s1(314);
  tmp_ivl_3059 <= state_in_s0(314);
  tmp_ivl_3060 <= tmp_ivl_3057 & tmp_ivl_3059;
  LPM_q_ivl_3063 <= tmp_ivl_3065 & tmp_ivl_3060;
  new_AGEMA_signal_2611 <= tmp_ivl_3069(1);
  tmp_ivl_3067 <= tmp_ivl_3069(0);
  tmp_ivl_3069 <= LPM_d0_ivl_3073(0 + 1 downto 0);
  tmp_ivl_3075 <= state_in_s1(293);
  tmp_ivl_3077 <= state_in_s0(293);
  tmp_ivl_3078 <= tmp_ivl_3075 & tmp_ivl_3077;
  LPM_q_ivl_3081 <= tmp_ivl_3083 & tmp_ivl_3078;
  tmp_ivl_3086 <= state_in_s1(37);
  tmp_ivl_3088 <= state_in_s0(37);
  tmp_ivl_3089 <= tmp_ivl_3086 & tmp_ivl_3088;
  LPM_q_ivl_3092 <= tmp_ivl_3094 & tmp_ivl_3089;
  new_AGEMA_signal_2613 <= tmp_ivl_3098(1);
  tmp_ivl_3096 <= tmp_ivl_3098(0);
  tmp_ivl_3098 <= LPM_d0_ivl_3102(0 + 1 downto 0);
  tmp_ivl_3104 <= state_in_s1(292);
  tmp_ivl_3106 <= state_in_s0(292);
  tmp_ivl_3107 <= tmp_ivl_3104 & tmp_ivl_3106;
  LPM_q_ivl_3110 <= tmp_ivl_3112 & tmp_ivl_3107;
  tmp_ivl_3115 <= state_in_s1(36);
  tmp_ivl_3117 <= state_in_s0(36);
  tmp_ivl_3118 <= tmp_ivl_3115 & tmp_ivl_3117;
  LPM_q_ivl_3121 <= tmp_ivl_3123 & tmp_ivl_3118;
  new_AGEMA_signal_2615 <= tmp_ivl_3127(1);
  tmp_ivl_3125 <= tmp_ivl_3127(0);
  tmp_ivl_3127 <= LPM_d0_ivl_3131(0 + 1 downto 0);
  tmp_ivl_3133 <= state_in_s1(35);
  tmp_ivl_3135 <= state_in_s0(35);
  tmp_ivl_3136 <= tmp_ivl_3133 & tmp_ivl_3135;
  LPM_q_ivl_3139 <= tmp_ivl_3141 & tmp_ivl_3136;
  tmp_ivl_3144 <= state_in_s1(291);
  tmp_ivl_3146 <= state_in_s0(291);
  tmp_ivl_3147 <= tmp_ivl_3144 & tmp_ivl_3146;
  LPM_q_ivl_3150 <= tmp_ivl_3152 & tmp_ivl_3147;
  new_AGEMA_signal_2617 <= tmp_ivl_3156(1);
  tmp_ivl_3154 <= tmp_ivl_3156(0);
  tmp_ivl_3156 <= LPM_d0_ivl_3160(0 + 1 downto 0);
  tmp_ivl_3162 <= state_in_s1(34);
  tmp_ivl_3164 <= state_in_s0(34);
  tmp_ivl_3165 <= tmp_ivl_3162 & tmp_ivl_3164;
  LPM_q_ivl_3168 <= tmp_ivl_3170 & tmp_ivl_3165;
  tmp_ivl_3173 <= state_in_s1(290);
  tmp_ivl_3175 <= state_in_s0(290);
  tmp_ivl_3176 <= tmp_ivl_3173 & tmp_ivl_3175;
  LPM_q_ivl_3179 <= tmp_ivl_3181 & tmp_ivl_3176;
  new_AGEMA_signal_2619 <= tmp_ivl_3185(1);
  tmp_ivl_3183 <= tmp_ivl_3185(0);
  tmp_ivl_3185 <= LPM_d0_ivl_3189(0 + 1 downto 0);
  tmp_ivl_3191 <= state_in_s1(289);
  tmp_ivl_3193 <= state_in_s0(289);
  tmp_ivl_3194 <= tmp_ivl_3191 & tmp_ivl_3193;
  LPM_q_ivl_3197 <= tmp_ivl_3199 & tmp_ivl_3194;
  tmp_ivl_3202 <= state_in_s1(33);
  tmp_ivl_3204 <= state_in_s0(33);
  tmp_ivl_3205 <= tmp_ivl_3202 & tmp_ivl_3204;
  LPM_q_ivl_3208 <= tmp_ivl_3210 & tmp_ivl_3205;
  new_AGEMA_signal_2621 <= tmp_ivl_3214(1);
  tmp_ivl_3212 <= tmp_ivl_3214(0);
  tmp_ivl_3214 <= LPM_d0_ivl_3218(0 + 1 downto 0);
  tmp_ivl_3220 <= state_in_s1(32);
  tmp_ivl_3222 <= state_in_s0(32);
  tmp_ivl_3223 <= tmp_ivl_3220 & tmp_ivl_3222;
  LPM_q_ivl_3226 <= tmp_ivl_3228 & tmp_ivl_3223;
  tmp_ivl_3231 <= state_in_s1(288);
  tmp_ivl_3233 <= state_in_s0(288);
  tmp_ivl_3234 <= tmp_ivl_3231 & tmp_ivl_3233;
  LPM_q_ivl_3237 <= tmp_ivl_3239 & tmp_ivl_3234;
  new_AGEMA_signal_2623 <= tmp_ivl_3243(1);
  tmp_ivl_3241 <= tmp_ivl_3243(0);
  tmp_ivl_3243 <= LPM_d0_ivl_3247(0 + 1 downto 0);
  tmp_ivl_3249 <= state_in_s1(47);
  tmp_ivl_3251 <= state_in_s0(47);
  tmp_ivl_3252 <= tmp_ivl_3249 & tmp_ivl_3251;
  LPM_q_ivl_3255 <= tmp_ivl_3257 & tmp_ivl_3252;
  tmp_ivl_3260 <= state_in_s1(303);
  tmp_ivl_3262 <= state_in_s0(303);
  tmp_ivl_3263 <= tmp_ivl_3260 & tmp_ivl_3262;
  LPM_q_ivl_3266 <= tmp_ivl_3268 & tmp_ivl_3263;
  new_AGEMA_signal_2625 <= tmp_ivl_3272(1);
  tmp_ivl_3270 <= tmp_ivl_3272(0);
  tmp_ivl_3272 <= LPM_d0_ivl_3276(0 + 1 downto 0);
  tmp_ivl_3278 <= state_in_s1(302);
  tmp_ivl_3280 <= state_in_s0(302);
  tmp_ivl_3281 <= tmp_ivl_3278 & tmp_ivl_3280;
  LPM_q_ivl_3284 <= tmp_ivl_3286 & tmp_ivl_3281;
  tmp_ivl_3289 <= state_in_s1(46);
  tmp_ivl_3291 <= state_in_s0(46);
  tmp_ivl_3292 <= tmp_ivl_3289 & tmp_ivl_3291;
  LPM_q_ivl_3295 <= tmp_ivl_3297 & tmp_ivl_3292;
  new_AGEMA_signal_2627 <= tmp_ivl_3301(1);
  tmp_ivl_3299 <= tmp_ivl_3301(0);
  tmp_ivl_3301 <= LPM_d0_ivl_3305(0 + 1 downto 0);
  tmp_ivl_3307 <= state_in_s1(45);
  tmp_ivl_3309 <= state_in_s0(45);
  tmp_ivl_3310 <= tmp_ivl_3307 & tmp_ivl_3309;
  LPM_q_ivl_3313 <= tmp_ivl_3315 & tmp_ivl_3310;
  tmp_ivl_3318 <= state_in_s1(301);
  tmp_ivl_3320 <= state_in_s0(301);
  tmp_ivl_3321 <= tmp_ivl_3318 & tmp_ivl_3320;
  LPM_q_ivl_3324 <= tmp_ivl_3326 & tmp_ivl_3321;
  new_AGEMA_signal_2629 <= tmp_ivl_3330(1);
  tmp_ivl_3328 <= tmp_ivl_3330(0);
  tmp_ivl_3330 <= LPM_d0_ivl_3334(0 + 1 downto 0);
  tmp_ivl_3336 <= state_in_s1(44);
  tmp_ivl_3338 <= state_in_s0(44);
  tmp_ivl_3339 <= tmp_ivl_3336 & tmp_ivl_3338;
  LPM_q_ivl_3342 <= tmp_ivl_3344 & tmp_ivl_3339;
  tmp_ivl_3347 <= state_in_s1(300);
  tmp_ivl_3349 <= state_in_s0(300);
  tmp_ivl_3350 <= tmp_ivl_3347 & tmp_ivl_3349;
  LPM_q_ivl_3353 <= tmp_ivl_3355 & tmp_ivl_3350;
  new_AGEMA_signal_2631 <= tmp_ivl_3359(1);
  tmp_ivl_3357 <= tmp_ivl_3359(0);
  tmp_ivl_3359 <= LPM_d0_ivl_3363(0 + 1 downto 0);
  tmp_ivl_3365 <= state_in_s1(57);
  tmp_ivl_3367 <= state_in_s0(57);
  tmp_ivl_3368 <= tmp_ivl_3365 & tmp_ivl_3367;
  LPM_q_ivl_3371 <= tmp_ivl_3373 & tmp_ivl_3368;
  tmp_ivl_3376 <= state_in_s1(313);
  tmp_ivl_3378 <= state_in_s0(313);
  tmp_ivl_3379 <= tmp_ivl_3376 & tmp_ivl_3378;
  LPM_q_ivl_3382 <= tmp_ivl_3384 & tmp_ivl_3379;
  new_AGEMA_signal_2633 <= tmp_ivl_3388(1);
  tmp_ivl_3386 <= tmp_ivl_3388(0);
  tmp_ivl_3388 <= LPM_d0_ivl_3392(0 + 1 downto 0);
  tmp_ivl_3394 <= state_in_s1(43);
  tmp_ivl_3396 <= state_in_s0(43);
  tmp_ivl_3397 <= tmp_ivl_3394 & tmp_ivl_3396;
  LPM_q_ivl_3400 <= tmp_ivl_3402 & tmp_ivl_3397;
  tmp_ivl_3405 <= state_in_s1(299);
  tmp_ivl_3407 <= state_in_s0(299);
  tmp_ivl_3408 <= tmp_ivl_3405 & tmp_ivl_3407;
  LPM_q_ivl_3411 <= tmp_ivl_3413 & tmp_ivl_3408;
  new_AGEMA_signal_2635 <= tmp_ivl_3417(1);
  tmp_ivl_3415 <= tmp_ivl_3417(0);
  tmp_ivl_3417 <= LPM_d0_ivl_3421(0 + 1 downto 0);
  tmp_ivl_3423 <= state_in_s1(298);
  tmp_ivl_3425 <= state_in_s0(298);
  tmp_ivl_3426 <= tmp_ivl_3423 & tmp_ivl_3425;
  LPM_q_ivl_3429 <= tmp_ivl_3431 & tmp_ivl_3426;
  tmp_ivl_3434 <= state_in_s1(42);
  tmp_ivl_3436 <= state_in_s0(42);
  tmp_ivl_3437 <= tmp_ivl_3434 & tmp_ivl_3436;
  LPM_q_ivl_3440 <= tmp_ivl_3442 & tmp_ivl_3437;
  new_AGEMA_signal_2637 <= tmp_ivl_3446(1);
  tmp_ivl_3444 <= tmp_ivl_3446(0);
  tmp_ivl_3446 <= LPM_d0_ivl_3450(0 + 1 downto 0);
  tmp_ivl_3452 <= state_in_s1(297);
  tmp_ivl_3454 <= state_in_s0(297);
  tmp_ivl_3455 <= tmp_ivl_3452 & tmp_ivl_3454;
  LPM_q_ivl_3458 <= tmp_ivl_3460 & tmp_ivl_3455;
  tmp_ivl_3463 <= state_in_s1(41);
  tmp_ivl_3465 <= state_in_s0(41);
  tmp_ivl_3466 <= tmp_ivl_3463 & tmp_ivl_3465;
  LPM_q_ivl_3469 <= tmp_ivl_3471 & tmp_ivl_3466;
  new_AGEMA_signal_2639 <= tmp_ivl_3475(1);
  tmp_ivl_3473 <= tmp_ivl_3475(0);
  tmp_ivl_3475 <= LPM_d0_ivl_3479(0 + 1 downto 0);
  tmp_ivl_3481 <= state_in_s1(40);
  tmp_ivl_3483 <= state_in_s0(40);
  tmp_ivl_3484 <= tmp_ivl_3481 & tmp_ivl_3483;
  LPM_q_ivl_3487 <= tmp_ivl_3489 & tmp_ivl_3484;
  tmp_ivl_3492 <= state_in_s1(296);
  tmp_ivl_3494 <= state_in_s0(296);
  tmp_ivl_3495 <= tmp_ivl_3492 & tmp_ivl_3494;
  LPM_q_ivl_3498 <= tmp_ivl_3500 & tmp_ivl_3495;
  new_AGEMA_signal_2641 <= tmp_ivl_3504(1);
  tmp_ivl_3502 <= tmp_ivl_3504(0);
  tmp_ivl_3504 <= LPM_d0_ivl_3508(0 + 1 downto 0);
  tmp_ivl_3510 <= state_in_s1(55);
  tmp_ivl_3512 <= state_in_s0(55);
  tmp_ivl_3513 <= tmp_ivl_3510 & tmp_ivl_3512;
  LPM_q_ivl_3516 <= tmp_ivl_3518 & tmp_ivl_3513;
  tmp_ivl_3521 <= state_in_s1(311);
  tmp_ivl_3523 <= state_in_s0(311);
  tmp_ivl_3524 <= tmp_ivl_3521 & tmp_ivl_3523;
  LPM_q_ivl_3527 <= tmp_ivl_3529 & tmp_ivl_3524;
  new_AGEMA_signal_2643 <= tmp_ivl_3533(1);
  tmp_ivl_3531 <= tmp_ivl_3533(0);
  tmp_ivl_3533 <= LPM_d0_ivl_3537(0 + 1 downto 0);
  tmp_ivl_3539 <= state_in_s1(54);
  tmp_ivl_3541 <= state_in_s0(54);
  tmp_ivl_3542 <= tmp_ivl_3539 & tmp_ivl_3541;
  LPM_q_ivl_3545 <= tmp_ivl_3547 & tmp_ivl_3542;
  tmp_ivl_3550 <= state_in_s1(310);
  tmp_ivl_3552 <= state_in_s0(310);
  tmp_ivl_3553 <= tmp_ivl_3550 & tmp_ivl_3552;
  LPM_q_ivl_3556 <= tmp_ivl_3558 & tmp_ivl_3553;
  new_AGEMA_signal_2645 <= tmp_ivl_3562(1);
  tmp_ivl_3560 <= tmp_ivl_3562(0);
  tmp_ivl_3562 <= LPM_d0_ivl_3566(0 + 1 downto 0);
  tmp_ivl_3568 <= state_in_s1(53);
  tmp_ivl_3570 <= state_in_s0(53);
  tmp_ivl_3571 <= tmp_ivl_3568 & tmp_ivl_3570;
  LPM_q_ivl_3574 <= tmp_ivl_3576 & tmp_ivl_3571;
  tmp_ivl_3579 <= state_in_s1(309);
  tmp_ivl_3581 <= state_in_s0(309);
  tmp_ivl_3582 <= tmp_ivl_3579 & tmp_ivl_3581;
  LPM_q_ivl_3585 <= tmp_ivl_3587 & tmp_ivl_3582;
  new_AGEMA_signal_2647 <= tmp_ivl_3591(1);
  tmp_ivl_3589 <= tmp_ivl_3591(0);
  tmp_ivl_3591 <= LPM_d0_ivl_3595(0 + 1 downto 0);
  tmp_ivl_3597 <= state_in_s1(52);
  tmp_ivl_3599 <= state_in_s0(52);
  tmp_ivl_3600 <= tmp_ivl_3597 & tmp_ivl_3599;
  LPM_q_ivl_3603 <= tmp_ivl_3605 & tmp_ivl_3600;
  tmp_ivl_3608 <= state_in_s1(308);
  tmp_ivl_3610 <= state_in_s0(308);
  tmp_ivl_3611 <= tmp_ivl_3608 & tmp_ivl_3610;
  LPM_q_ivl_3614 <= tmp_ivl_3616 & tmp_ivl_3611;
  new_AGEMA_signal_2649 <= tmp_ivl_3620(1);
  tmp_ivl_3618 <= tmp_ivl_3620(0);
  tmp_ivl_3620 <= LPM_d0_ivl_3624(0 + 1 downto 0);
  tmp_ivl_3626 <= state_in_s1(307);
  tmp_ivl_3628 <= state_in_s0(307);
  tmp_ivl_3629 <= tmp_ivl_3626 & tmp_ivl_3628;
  LPM_q_ivl_3632 <= tmp_ivl_3634 & tmp_ivl_3629;
  tmp_ivl_3637 <= state_in_s1(51);
  tmp_ivl_3639 <= state_in_s0(51);
  tmp_ivl_3640 <= tmp_ivl_3637 & tmp_ivl_3639;
  LPM_q_ivl_3643 <= tmp_ivl_3645 & tmp_ivl_3640;
  new_AGEMA_signal_2651 <= tmp_ivl_3649(1);
  tmp_ivl_3647 <= tmp_ivl_3649(0);
  tmp_ivl_3649 <= LPM_d0_ivl_3653(0 + 1 downto 0);
  tmp_ivl_3655 <= state_in_s1(50);
  tmp_ivl_3657 <= state_in_s0(50);
  tmp_ivl_3658 <= tmp_ivl_3655 & tmp_ivl_3657;
  LPM_q_ivl_3661 <= tmp_ivl_3663 & tmp_ivl_3658;
  tmp_ivl_3666 <= state_in_s1(306);
  tmp_ivl_3668 <= state_in_s0(306);
  tmp_ivl_3669 <= tmp_ivl_3666 & tmp_ivl_3668;
  LPM_q_ivl_3672 <= tmp_ivl_3674 & tmp_ivl_3669;
  new_AGEMA_signal_2653 <= tmp_ivl_3678(1);
  tmp_ivl_3676 <= tmp_ivl_3678(0);
  tmp_ivl_3678 <= LPM_d0_ivl_3682(0 + 1 downto 0);
  tmp_ivl_3684 <= state_in_s1(56);
  tmp_ivl_3686 <= state_in_s0(56);
  tmp_ivl_3687 <= tmp_ivl_3684 & tmp_ivl_3686;
  LPM_q_ivl_3690 <= tmp_ivl_3692 & tmp_ivl_3687;
  tmp_ivl_3695 <= state_in_s1(312);
  tmp_ivl_3697 <= state_in_s0(312);
  tmp_ivl_3698 <= tmp_ivl_3695 & tmp_ivl_3697;
  LPM_q_ivl_3701 <= tmp_ivl_3703 & tmp_ivl_3698;
  new_AGEMA_signal_2655 <= tmp_ivl_3707(1);
  tmp_ivl_3705 <= tmp_ivl_3707(0);
  tmp_ivl_3707 <= LPM_d0_ivl_3711(0 + 1 downto 0);
  tmp_ivl_3713 <= state_in_s1(66);
  tmp_ivl_3715 <= state_in_s0(66);
  tmp_ivl_3716 <= tmp_ivl_3713 & tmp_ivl_3715;
  LPM_q_ivl_3719 <= tmp_ivl_3721 & tmp_ivl_3716;
  tmp_ivl_3724 <= state_in_s1(258);
  tmp_ivl_3726 <= state_in_s0(258);
  tmp_ivl_3727 <= tmp_ivl_3724 & tmp_ivl_3726;
  LPM_q_ivl_3730 <= tmp_ivl_3732 & tmp_ivl_3727;
  new_AGEMA_signal_2657 <= tmp_ivl_3734(1);
  n3310 <= tmp_ivl_3734(0);
  tmp_ivl_3734 <= LPM_d0_ivl_3738(0 + 1 downto 0);
  tmp_ivl_3740 <= state_in_s1(67);
  tmp_ivl_3742 <= state_in_s0(67);
  tmp_ivl_3743 <= tmp_ivl_3740 & tmp_ivl_3742;
  LPM_q_ivl_3746 <= tmp_ivl_3748 & tmp_ivl_3743;
  tmp_ivl_3751 <= state_in_s1(259);
  tmp_ivl_3753 <= state_in_s0(259);
  tmp_ivl_3754 <= tmp_ivl_3751 & tmp_ivl_3753;
  LPM_q_ivl_3757 <= tmp_ivl_3759 & tmp_ivl_3754;
  new_AGEMA_signal_2659 <= tmp_ivl_3761(1);
  n3317 <= tmp_ivl_3761(0);
  tmp_ivl_3761 <= LPM_d0_ivl_3765(0 + 1 downto 0);
  tmp_ivl_3767 <= state_in_s1(65);
  tmp_ivl_3769 <= state_in_s0(65);
  tmp_ivl_3770 <= tmp_ivl_3767 & tmp_ivl_3769;
  LPM_q_ivl_3773 <= tmp_ivl_3775 & tmp_ivl_3770;
  tmp_ivl_3778 <= state_in_s1(257);
  tmp_ivl_3780 <= state_in_s0(257);
  tmp_ivl_3781 <= tmp_ivl_3778 & tmp_ivl_3780;
  LPM_q_ivl_3784 <= tmp_ivl_3786 & tmp_ivl_3781;
  new_AGEMA_signal_2661 <= tmp_ivl_3788(1);
  n3329 <= tmp_ivl_3788(0);
  tmp_ivl_3788 <= LPM_d0_ivl_3792(0 + 1 downto 0);
  tmp_ivl_3794 <= state_in_s1(106);
  tmp_ivl_3796 <= state_in_s0(106);
  tmp_ivl_3797 <= tmp_ivl_3794 & tmp_ivl_3796;
  LPM_q_ivl_3800 <= tmp_ivl_3802 & tmp_ivl_3797;
  tmp_ivl_3805 <= state_in_s1(298);
  tmp_ivl_3807 <= state_in_s0(298);
  tmp_ivl_3808 <= tmp_ivl_3805 & tmp_ivl_3807;
  LPM_q_ivl_3811 <= tmp_ivl_3813 & tmp_ivl_3808;
  new_AGEMA_signal_2663 <= tmp_ivl_3815(1);
  n3336 <= tmp_ivl_3815(0);
  tmp_ivl_3815 <= LPM_d0_ivl_3819(0 + 1 downto 0);
  tmp_ivl_3821 <= state_in_s1(105);
  tmp_ivl_3823 <= state_in_s0(105);
  tmp_ivl_3824 <= tmp_ivl_3821 & tmp_ivl_3823;
  LPM_q_ivl_3827 <= tmp_ivl_3829 & tmp_ivl_3824;
  tmp_ivl_3832 <= state_in_s1(297);
  tmp_ivl_3834 <= state_in_s0(297);
  tmp_ivl_3835 <= tmp_ivl_3832 & tmp_ivl_3834;
  LPM_q_ivl_3838 <= tmp_ivl_3840 & tmp_ivl_3835;
  new_AGEMA_signal_2665 <= tmp_ivl_3842(1);
  n3348 <= tmp_ivl_3842(0);
  tmp_ivl_3842 <= LPM_d0_ivl_3846(0 + 1 downto 0);
  tmp_ivl_3848 <= state_in_s1(97);
  tmp_ivl_3850 <= state_in_s0(97);
  tmp_ivl_3851 <= tmp_ivl_3848 & tmp_ivl_3850;
  LPM_q_ivl_3854 <= tmp_ivl_3856 & tmp_ivl_3851;
  tmp_ivl_3859 <= state_in_s1(289);
  tmp_ivl_3861 <= state_in_s0(289);
  tmp_ivl_3862 <= tmp_ivl_3859 & tmp_ivl_3861;
  LPM_q_ivl_3865 <= tmp_ivl_3867 & tmp_ivl_3862;
  new_AGEMA_signal_2667 <= tmp_ivl_3869(1);
  n3367 <= tmp_ivl_3869(0);
  tmp_ivl_3869 <= LPM_d0_ivl_3873(0 + 1 downto 0);
  tmp_ivl_3875 <= state_in_s1(87);
  tmp_ivl_3877 <= state_in_s0(87);
  tmp_ivl_3878 <= tmp_ivl_3875 & tmp_ivl_3877;
  LPM_q_ivl_3881 <= tmp_ivl_3883 & tmp_ivl_3878;
  tmp_ivl_3886 <= state_in_s1(279);
  tmp_ivl_3888 <= state_in_s0(279);
  tmp_ivl_3889 <= tmp_ivl_3886 & tmp_ivl_3888;
  LPM_q_ivl_3892 <= tmp_ivl_3894 & tmp_ivl_3889;
  new_AGEMA_signal_2669 <= tmp_ivl_3896(1);
  n3370 <= tmp_ivl_3896(0);
  tmp_ivl_3896 <= LPM_d0_ivl_3900(0 + 1 downto 0);
  tmp_ivl_3902 <= state_in_s1(72);
  tmp_ivl_3904 <= state_in_s0(72);
  tmp_ivl_3905 <= tmp_ivl_3902 & tmp_ivl_3904;
  LPM_q_ivl_3908 <= tmp_ivl_3910 & tmp_ivl_3905;
  tmp_ivl_3913 <= state_in_s1(264);
  tmp_ivl_3915 <= state_in_s0(264);
  tmp_ivl_3916 <= tmp_ivl_3913 & tmp_ivl_3915;
  LPM_q_ivl_3919 <= tmp_ivl_3921 & tmp_ivl_3916;
  new_AGEMA_signal_2671 <= tmp_ivl_3923(1);
  n3386 <= tmp_ivl_3923(0);
  tmp_ivl_3923 <= LPM_d0_ivl_3927(0 + 1 downto 0);
  tmp_ivl_3929 <= state_in_s1(75);
  tmp_ivl_3931 <= state_in_s0(75);
  tmp_ivl_3932 <= tmp_ivl_3929 & tmp_ivl_3931;
  LPM_q_ivl_3935 <= tmp_ivl_3937 & tmp_ivl_3932;
  tmp_ivl_3940 <= state_in_s1(267);
  tmp_ivl_3942 <= state_in_s0(267);
  tmp_ivl_3943 <= tmp_ivl_3940 & tmp_ivl_3942;
  LPM_q_ivl_3946 <= tmp_ivl_3948 & tmp_ivl_3943;
  new_AGEMA_signal_2673 <= tmp_ivl_3950(1);
  n3388 <= tmp_ivl_3950(0);
  tmp_ivl_3950 <= LPM_d0_ivl_3954(0 + 1 downto 0);
  tmp_ivl_3956 <= state_in_s1(76);
  tmp_ivl_3958 <= state_in_s0(76);
  tmp_ivl_3959 <= tmp_ivl_3956 & tmp_ivl_3958;
  LPM_q_ivl_3962 <= tmp_ivl_3964 & tmp_ivl_3959;
  tmp_ivl_3967 <= state_in_s1(268);
  tmp_ivl_3969 <= state_in_s0(268);
  tmp_ivl_3970 <= tmp_ivl_3967 & tmp_ivl_3969;
  LPM_q_ivl_3973 <= tmp_ivl_3975 & tmp_ivl_3970;
  new_AGEMA_signal_2675 <= tmp_ivl_3977(1);
  n3430 <= tmp_ivl_3977(0);
  tmp_ivl_3977 <= LPM_d0_ivl_3981(0 + 1 downto 0);
  tmp_ivl_3983 <= state_in_s1(115);
  tmp_ivl_3985 <= state_in_s0(115);
  tmp_ivl_3986 <= tmp_ivl_3983 & tmp_ivl_3985;
  LPM_q_ivl_3989 <= tmp_ivl_3991 & tmp_ivl_3986;
  tmp_ivl_3994 <= state_in_s1(307);
  tmp_ivl_3996 <= state_in_s0(307);
  tmp_ivl_3997 <= tmp_ivl_3994 & tmp_ivl_3996;
  LPM_q_ivl_4000 <= tmp_ivl_4002 & tmp_ivl_3997;
  new_AGEMA_signal_2677 <= tmp_ivl_4004(1);
  n3449 <= tmp_ivl_4004(0);
  tmp_ivl_4004 <= LPM_d0_ivl_4008(0 + 1 downto 0);
  tmp_ivl_4010 <= state_in_s1(100);
  tmp_ivl_4012 <= state_in_s0(100);
  tmp_ivl_4013 <= tmp_ivl_4010 & tmp_ivl_4012;
  LPM_q_ivl_4016 <= tmp_ivl_4018 & tmp_ivl_4013;
  tmp_ivl_4021 <= state_in_s1(292);
  tmp_ivl_4023 <= state_in_s0(292);
  tmp_ivl_4024 <= tmp_ivl_4021 & tmp_ivl_4023;
  LPM_q_ivl_4027 <= tmp_ivl_4029 & tmp_ivl_4024;
  new_AGEMA_signal_2679 <= tmp_ivl_4031(1);
  n3469 <= tmp_ivl_4031(0);
  tmp_ivl_4031 <= LPM_d0_ivl_4035(0 + 1 downto 0);
  tmp_ivl_4037 <= state_in_s1(101);
  tmp_ivl_4039 <= state_in_s0(101);
  tmp_ivl_4040 <= tmp_ivl_4037 & tmp_ivl_4039;
  LPM_q_ivl_4043 <= tmp_ivl_4045 & tmp_ivl_4040;
  tmp_ivl_4048 <= state_in_s1(293);
  tmp_ivl_4050 <= state_in_s0(293);
  tmp_ivl_4051 <= tmp_ivl_4048 & tmp_ivl_4050;
  LPM_q_ivl_4054 <= tmp_ivl_4056 & tmp_ivl_4051;
  new_AGEMA_signal_2681 <= tmp_ivl_4058(1);
  n3520 <= tmp_ivl_4058(0);
  tmp_ivl_4058 <= LPM_d0_ivl_4062(0 + 1 downto 0);
  tmp_ivl_4064 <= state_in_s1(110);
  tmp_ivl_4066 <= state_in_s0(110);
  tmp_ivl_4067 <= tmp_ivl_4064 & tmp_ivl_4066;
  LPM_q_ivl_4070 <= tmp_ivl_4072 & tmp_ivl_4067;
  tmp_ivl_4075 <= state_in_s1(302);
  tmp_ivl_4077 <= state_in_s0(302);
  tmp_ivl_4078 <= tmp_ivl_4075 & tmp_ivl_4077;
  LPM_q_ivl_4081 <= tmp_ivl_4083 & tmp_ivl_4078;
  new_AGEMA_signal_2683 <= tmp_ivl_4085(1);
  n3547 <= tmp_ivl_4085(0);
  tmp_ivl_4085 <= LPM_d0_ivl_4089(0 + 1 downto 0);
  tmp_ivl_4091 <= state_in_s1(81);
  tmp_ivl_4093 <= state_in_s0(81);
  tmp_ivl_4094 <= tmp_ivl_4091 & tmp_ivl_4093;
  LPM_q_ivl_4097 <= tmp_ivl_4099 & tmp_ivl_4094;
  tmp_ivl_4102 <= state_in_s1(273);
  tmp_ivl_4104 <= state_in_s0(273);
  tmp_ivl_4105 <= tmp_ivl_4102 & tmp_ivl_4104;
  LPM_q_ivl_4108 <= tmp_ivl_4110 & tmp_ivl_4105;
  new_AGEMA_signal_2685 <= tmp_ivl_4112(1);
  n3610 <= tmp_ivl_4112(0);
  tmp_ivl_4112 <= LPM_d0_ivl_4116(0 + 1 downto 0);
  tmp_ivl_4118 <= state_in_s1(84);
  tmp_ivl_4120 <= state_in_s0(84);
  tmp_ivl_4121 <= tmp_ivl_4118 & tmp_ivl_4120;
  LPM_q_ivl_4124 <= tmp_ivl_4126 & tmp_ivl_4121;
  tmp_ivl_4129 <= state_in_s1(276);
  tmp_ivl_4131 <= state_in_s0(276);
  tmp_ivl_4132 <= tmp_ivl_4129 & tmp_ivl_4131;
  LPM_q_ivl_4135 <= tmp_ivl_4137 & tmp_ivl_4132;
  new_AGEMA_signal_2687 <= tmp_ivl_4139(1);
  n3699 <= tmp_ivl_4139(0);
  tmp_ivl_4139 <= LPM_d0_ivl_4143(0 + 1 downto 0);
  tmp_ivl_4145 <= state_in_s1(85);
  tmp_ivl_4147 <= state_in_s0(85);
  tmp_ivl_4148 <= tmp_ivl_4145 & tmp_ivl_4147;
  LPM_q_ivl_4151 <= tmp_ivl_4153 & tmp_ivl_4148;
  tmp_ivl_4156 <= state_in_s1(277);
  tmp_ivl_4158 <= state_in_s0(277);
  tmp_ivl_4159 <= tmp_ivl_4156 & tmp_ivl_4158;
  LPM_q_ivl_4162 <= tmp_ivl_4164 & tmp_ivl_4159;
  new_AGEMA_signal_2689 <= tmp_ivl_4166(1);
  n3793 <= tmp_ivl_4166(0);
  tmp_ivl_4166 <= LPM_d0_ivl_4170(0 + 1 downto 0);
  tmp_ivl_4172 <= state_in_s1(177);
  tmp_ivl_4174 <= state_in_s0(177);
  tmp_ivl_4175 <= tmp_ivl_4172 & tmp_ivl_4174;
  LPM_q_ivl_4178 <= tmp_ivl_4180 & tmp_ivl_4175;
  tmp_ivl_4183 <= state_in_s1(113);
  tmp_ivl_4185 <= state_in_s0(113);
  tmp_ivl_4186 <= tmp_ivl_4183 & tmp_ivl_4185;
  LPM_q_ivl_4189 <= tmp_ivl_4191 & tmp_ivl_4186;
  new_AGEMA_signal_2692 <= tmp_ivl_4193(1);
  n3291 <= tmp_ivl_4193(0);
  tmp_ivl_4193 <= LPM_d0_ivl_4197(0 + 1 downto 0);
  tmp_ivl_4199 <= state_in_s1(171);
  tmp_ivl_4201 <= state_in_s0(171);
  tmp_ivl_4202 <= tmp_ivl_4199 & tmp_ivl_4201;
  LPM_q_ivl_4205 <= tmp_ivl_4207 & tmp_ivl_4202;
  tmp_ivl_4210 <= state_in_s1(107);
  tmp_ivl_4212 <= state_in_s0(107);
  tmp_ivl_4213 <= tmp_ivl_4210 & tmp_ivl_4212;
  LPM_q_ivl_4216 <= tmp_ivl_4218 & tmp_ivl_4213;
  new_AGEMA_signal_2695 <= tmp_ivl_4220(1);
  n3280 <= tmp_ivl_4220(0);
  tmp_ivl_4220 <= LPM_d0_ivl_4224(0 + 1 downto 0);
  tmp_ivl_4226 <= state_in_s1(98);
  tmp_ivl_4228 <= state_in_s0(98);
  tmp_ivl_4229 <= tmp_ivl_4226 & tmp_ivl_4228;
  LPM_q_ivl_4232 <= tmp_ivl_4234 & tmp_ivl_4229;
  tmp_ivl_4237 <= state_in_s1(162);
  tmp_ivl_4239 <= state_in_s0(162);
  tmp_ivl_4240 <= tmp_ivl_4237 & tmp_ivl_4239;
  LPM_q_ivl_4243 <= tmp_ivl_4245 & tmp_ivl_4240;
  new_AGEMA_signal_2698 <= tmp_ivl_4247(1);
  n3273 <= tmp_ivl_4247(0);
  tmp_ivl_4247 <= LPM_d0_ivl_4251(0 + 1 downto 0);
  tmp_ivl_4253 <= state_in_s1(172);
  tmp_ivl_4255 <= state_in_s0(172);
  tmp_ivl_4256 <= tmp_ivl_4253 & tmp_ivl_4255;
  LPM_q_ivl_4259 <= tmp_ivl_4261 & tmp_ivl_4256;
  tmp_ivl_4264 <= state_in_s1(108);
  tmp_ivl_4266 <= state_in_s0(108);
  tmp_ivl_4267 <= tmp_ivl_4264 & tmp_ivl_4266;
  LPM_q_ivl_4270 <= tmp_ivl_4272 & tmp_ivl_4267;
  new_AGEMA_signal_2701 <= tmp_ivl_4274(1);
  n3279 <= tmp_ivl_4274(0);
  tmp_ivl_4274 <= LPM_d0_ivl_4278(0 + 1 downto 0);
  tmp_ivl_4280 <= state_in_s1(178);
  tmp_ivl_4282 <= state_in_s0(178);
  tmp_ivl_4283 <= tmp_ivl_4280 & tmp_ivl_4282;
  LPM_q_ivl_4286 <= tmp_ivl_4288 & tmp_ivl_4283;
  tmp_ivl_4291 <= state_in_s1(114);
  tmp_ivl_4293 <= state_in_s0(114);
  tmp_ivl_4294 <= tmp_ivl_4291 & tmp_ivl_4293;
  LPM_q_ivl_4297 <= tmp_ivl_4299 & tmp_ivl_4294;
  new_AGEMA_signal_2704 <= tmp_ivl_4301(1);
  n3290 <= tmp_ivl_4301(0);
  tmp_ivl_4301 <= LPM_d0_ivl_4305(0 + 1 downto 0);
  tmp_ivl_4307 <= state_in_s1(99);
  tmp_ivl_4309 <= state_in_s0(99);
  tmp_ivl_4310 <= tmp_ivl_4307 & tmp_ivl_4309;
  LPM_q_ivl_4313 <= tmp_ivl_4315 & tmp_ivl_4310;
  tmp_ivl_4318 <= state_in_s1(163);
  tmp_ivl_4320 <= state_in_s0(163);
  tmp_ivl_4321 <= tmp_ivl_4318 & tmp_ivl_4320;
  LPM_q_ivl_4324 <= tmp_ivl_4326 & tmp_ivl_4321;
  new_AGEMA_signal_2707 <= tmp_ivl_4328(1);
  n3272 <= tmp_ivl_4328(0);
  tmp_ivl_4328 <= LPM_d0_ivl_4332(0 + 1 downto 0);
  tmp_ivl_4334 <= state_in_s1(115);
  tmp_ivl_4336 <= state_in_s0(115);
  tmp_ivl_4337 <= tmp_ivl_4334 & tmp_ivl_4336;
  LPM_q_ivl_4340 <= tmp_ivl_4342 & tmp_ivl_4337;
  tmp_ivl_4345 <= state_in_s1(179);
  tmp_ivl_4347 <= state_in_s0(179);
  tmp_ivl_4348 <= tmp_ivl_4345 & tmp_ivl_4347;
  LPM_q_ivl_4351 <= tmp_ivl_4353 & tmp_ivl_4348;
  new_AGEMA_signal_2709 <= tmp_ivl_4355(1);
  n3289 <= tmp_ivl_4355(0);
  tmp_ivl_4355 <= LPM_d0_ivl_4359(0 + 1 downto 0);
  tmp_ivl_4361 <= state_in_s1(109);
  tmp_ivl_4363 <= state_in_s0(109);
  tmp_ivl_4364 <= tmp_ivl_4361 & tmp_ivl_4363;
  LPM_q_ivl_4367 <= tmp_ivl_4369 & tmp_ivl_4364;
  tmp_ivl_4372 <= state_in_s1(173);
  tmp_ivl_4374 <= state_in_s0(173);
  tmp_ivl_4375 <= tmp_ivl_4372 & tmp_ivl_4374;
  LPM_q_ivl_4378 <= tmp_ivl_4380 & tmp_ivl_4375;
  new_AGEMA_signal_2712 <= tmp_ivl_4382(1);
  n3278 <= tmp_ivl_4382(0);
  tmp_ivl_4382 <= LPM_d0_ivl_4386(0 + 1 downto 0);
  tmp_ivl_4388 <= state_in_s1(100);
  tmp_ivl_4390 <= state_in_s0(100);
  tmp_ivl_4391 <= tmp_ivl_4388 & tmp_ivl_4390;
  LPM_q_ivl_4394 <= tmp_ivl_4396 & tmp_ivl_4391;
  tmp_ivl_4399 <= state_in_s1(164);
  tmp_ivl_4401 <= state_in_s0(164);
  tmp_ivl_4402 <= tmp_ivl_4399 & tmp_ivl_4401;
  LPM_q_ivl_4405 <= tmp_ivl_4407 & tmp_ivl_4402;
  new_AGEMA_signal_2714 <= tmp_ivl_4409(1);
  n3271 <= tmp_ivl_4409(0);
  tmp_ivl_4409 <= LPM_d0_ivl_4413(0 + 1 downto 0);
  tmp_ivl_4415 <= state_in_s1(180);
  tmp_ivl_4417 <= state_in_s0(180);
  tmp_ivl_4418 <= tmp_ivl_4415 & tmp_ivl_4417;
  LPM_q_ivl_4421 <= tmp_ivl_4423 & tmp_ivl_4418;
  tmp_ivl_4426 <= state_in_s1(116);
  tmp_ivl_4428 <= state_in_s0(116);
  tmp_ivl_4429 <= tmp_ivl_4426 & tmp_ivl_4428;
  LPM_q_ivl_4432 <= tmp_ivl_4434 & tmp_ivl_4429;
  new_AGEMA_signal_2717 <= tmp_ivl_4436(1);
  n3288 <= tmp_ivl_4436(0);
  tmp_ivl_4436 <= LPM_d0_ivl_4440(0 + 1 downto 0);
  tmp_ivl_4442 <= state_in_s1(110);
  tmp_ivl_4444 <= state_in_s0(110);
  tmp_ivl_4445 <= tmp_ivl_4442 & tmp_ivl_4444;
  LPM_q_ivl_4448 <= tmp_ivl_4450 & tmp_ivl_4445;
  tmp_ivl_4453 <= state_in_s1(174);
  tmp_ivl_4455 <= state_in_s0(174);
  tmp_ivl_4456 <= tmp_ivl_4453 & tmp_ivl_4455;
  LPM_q_ivl_4459 <= tmp_ivl_4461 & tmp_ivl_4456;
  new_AGEMA_signal_2719 <= tmp_ivl_4463(1);
  n3277 <= tmp_ivl_4463(0);
  tmp_ivl_4463 <= LPM_d0_ivl_4467(0 + 1 downto 0);
  tmp_ivl_4469 <= state_in_s1(101);
  tmp_ivl_4471 <= state_in_s0(101);
  tmp_ivl_4472 <= tmp_ivl_4469 & tmp_ivl_4471;
  LPM_q_ivl_4475 <= tmp_ivl_4477 & tmp_ivl_4472;
  tmp_ivl_4480 <= state_in_s1(165);
  tmp_ivl_4482 <= state_in_s0(165);
  tmp_ivl_4483 <= tmp_ivl_4480 & tmp_ivl_4482;
  LPM_q_ivl_4486 <= tmp_ivl_4488 & tmp_ivl_4483;
  new_AGEMA_signal_2721 <= tmp_ivl_4490(1);
  n3270 <= tmp_ivl_4490(0);
  tmp_ivl_4490 <= LPM_d0_ivl_4494(0 + 1 downto 0);
  tmp_ivl_4496 <= state_in_s1(175);
  tmp_ivl_4498 <= state_in_s0(175);
  tmp_ivl_4499 <= tmp_ivl_4496 & tmp_ivl_4498;
  LPM_q_ivl_4502 <= tmp_ivl_4504 & tmp_ivl_4499;
  tmp_ivl_4507 <= state_in_s1(111);
  tmp_ivl_4509 <= state_in_s0(111);
  tmp_ivl_4510 <= tmp_ivl_4507 & tmp_ivl_4509;
  LPM_q_ivl_4513 <= tmp_ivl_4515 & tmp_ivl_4510;
  new_AGEMA_signal_2724 <= tmp_ivl_4517(1);
  n3276 <= tmp_ivl_4517(0);
  tmp_ivl_4517 <= LPM_d0_ivl_4521(0 + 1 downto 0);
  tmp_ivl_4523 <= state_in_s1(181);
  tmp_ivl_4525 <= state_in_s0(181);
  tmp_ivl_4526 <= tmp_ivl_4523 & tmp_ivl_4525;
  LPM_q_ivl_4529 <= tmp_ivl_4531 & tmp_ivl_4526;
  tmp_ivl_4534 <= state_in_s1(117);
  tmp_ivl_4536 <= state_in_s0(117);
  tmp_ivl_4537 <= tmp_ivl_4534 & tmp_ivl_4536;
  LPM_q_ivl_4540 <= tmp_ivl_4542 & tmp_ivl_4537;
  new_AGEMA_signal_2727 <= tmp_ivl_4544(1);
  n3286 <= tmp_ivl_4544(0);
  tmp_ivl_4544 <= LPM_d0_ivl_4548(0 + 1 downto 0);
  tmp_ivl_4550 <= state_in_s1(102);
  tmp_ivl_4552 <= state_in_s0(102);
  tmp_ivl_4553 <= tmp_ivl_4550 & tmp_ivl_4552;
  LPM_q_ivl_4556 <= tmp_ivl_4558 & tmp_ivl_4553;
  tmp_ivl_4561 <= state_in_s1(166);
  tmp_ivl_4563 <= state_in_s0(166);
  tmp_ivl_4564 <= tmp_ivl_4561 & tmp_ivl_4563;
  LPM_q_ivl_4567 <= tmp_ivl_4569 & tmp_ivl_4564;
  new_AGEMA_signal_2730 <= tmp_ivl_4571(1);
  n3269 <= tmp_ivl_4571(0);
  tmp_ivl_4571 <= LPM_d0_ivl_4575(0 + 1 downto 0);
  tmp_ivl_4577 <= state_in_s1(182);
  tmp_ivl_4579 <= state_in_s0(182);
  tmp_ivl_4580 <= tmp_ivl_4577 & tmp_ivl_4579;
  LPM_q_ivl_4583 <= tmp_ivl_4585 & tmp_ivl_4580;
  tmp_ivl_4588 <= state_in_s1(118);
  tmp_ivl_4590 <= state_in_s0(118);
  tmp_ivl_4591 <= tmp_ivl_4588 & tmp_ivl_4590;
  LPM_q_ivl_4594 <= tmp_ivl_4596 & tmp_ivl_4591;
  new_AGEMA_signal_2733 <= tmp_ivl_4598(1);
  n3285 <= tmp_ivl_4598(0);
  tmp_ivl_4598 <= LPM_d0_ivl_4602(0 + 1 downto 0);
  tmp_ivl_4604 <= state_in_s1(160);
  tmp_ivl_4606 <= state_in_s0(160);
  tmp_ivl_4607 <= tmp_ivl_4604 & tmp_ivl_4606;
  LPM_q_ivl_4610 <= tmp_ivl_4612 & tmp_ivl_4607;
  tmp_ivl_4615 <= state_in_s1(96);
  tmp_ivl_4617 <= state_in_s0(96);
  tmp_ivl_4618 <= tmp_ivl_4615 & tmp_ivl_4617;
  LPM_q_ivl_4621 <= tmp_ivl_4623 & tmp_ivl_4618;
  new_AGEMA_signal_2736 <= tmp_ivl_4625(1);
  n3275 <= tmp_ivl_4625(0);
  tmp_ivl_4625 <= LPM_d0_ivl_4629(0 + 1 downto 0);
  tmp_ivl_4631 <= state_in_s1(103);
  tmp_ivl_4633 <= state_in_s0(103);
  tmp_ivl_4634 <= tmp_ivl_4631 & tmp_ivl_4633;
  LPM_q_ivl_4637 <= tmp_ivl_4639 & tmp_ivl_4634;
  tmp_ivl_4642 <= state_in_s1(167);
  tmp_ivl_4644 <= state_in_s0(167);
  tmp_ivl_4645 <= tmp_ivl_4642 & tmp_ivl_4644;
  LPM_q_ivl_4648 <= tmp_ivl_4650 & tmp_ivl_4645;
  new_AGEMA_signal_2739 <= tmp_ivl_4652(1);
  n3268 <= tmp_ivl_4652(0);
  tmp_ivl_4652 <= LPM_d0_ivl_4656(0 + 1 downto 0);
  tmp_ivl_4658 <= state_in_s1(119);
  tmp_ivl_4660 <= state_in_s0(119);
  tmp_ivl_4661 <= tmp_ivl_4658 & tmp_ivl_4660;
  LPM_q_ivl_4664 <= tmp_ivl_4666 & tmp_ivl_4661;
  tmp_ivl_4669 <= state_in_s1(183);
  tmp_ivl_4671 <= state_in_s0(183);
  tmp_ivl_4672 <= tmp_ivl_4669 & tmp_ivl_4671;
  LPM_q_ivl_4675 <= tmp_ivl_4677 & tmp_ivl_4672;
  new_AGEMA_signal_2742 <= tmp_ivl_4679(1);
  n3284 <= tmp_ivl_4679(0);
  tmp_ivl_4679 <= LPM_d0_ivl_4683(0 + 1 downto 0);
  tmp_ivl_4685 <= state_in_s1(97);
  tmp_ivl_4687 <= state_in_s0(97);
  tmp_ivl_4688 <= tmp_ivl_4685 & tmp_ivl_4687;
  LPM_q_ivl_4691 <= tmp_ivl_4693 & tmp_ivl_4688;
  tmp_ivl_4696 <= state_in_s1(161);
  tmp_ivl_4698 <= state_in_s0(161);
  tmp_ivl_4699 <= tmp_ivl_4696 & tmp_ivl_4698;
  LPM_q_ivl_4702 <= tmp_ivl_4704 & tmp_ivl_4699;
  new_AGEMA_signal_2744 <= tmp_ivl_4706(1);
  n3274 <= tmp_ivl_4706(0);
  tmp_ivl_4706 <= LPM_d0_ivl_4710(0 + 1 downto 0);
  tmp_ivl_4712 <= state_in_s1(88);
  tmp_ivl_4714 <= state_in_s0(88);
  tmp_ivl_4715 <= tmp_ivl_4712 & tmp_ivl_4714;
  LPM_q_ivl_4718 <= tmp_ivl_4720 & tmp_ivl_4715;
  tmp_ivl_4723 <= state_in_s1(152);
  tmp_ivl_4725 <= state_in_s0(152);
  tmp_ivl_4726 <= tmp_ivl_4723 & tmp_ivl_4725;
  LPM_q_ivl_4729 <= tmp_ivl_4731 & tmp_ivl_4726;
  new_AGEMA_signal_2747 <= tmp_ivl_4733(1);
  n3267 <= tmp_ivl_4733(0);
  tmp_ivl_4733 <= LPM_d0_ivl_4737(0 + 1 downto 0);
  tmp_ivl_4739 <= state_in_s1(168);
  tmp_ivl_4741 <= state_in_s0(168);
  tmp_ivl_4742 <= tmp_ivl_4739 & tmp_ivl_4741;
  LPM_q_ivl_4745 <= tmp_ivl_4747 & tmp_ivl_4742;
  tmp_ivl_4750 <= state_in_s1(104);
  tmp_ivl_4752 <= state_in_s0(104);
  tmp_ivl_4753 <= tmp_ivl_4750 & tmp_ivl_4752;
  LPM_q_ivl_4756 <= tmp_ivl_4758 & tmp_ivl_4753;
  new_AGEMA_signal_2750 <= tmp_ivl_4760(1);
  n3283 <= tmp_ivl_4760(0);
  tmp_ivl_4760 <= LPM_d0_ivl_4764(0 + 1 downto 0);
  tmp_ivl_4766 <= state_in_s1(89);
  tmp_ivl_4768 <= state_in_s0(89);
  tmp_ivl_4769 <= tmp_ivl_4766 & tmp_ivl_4768;
  LPM_q_ivl_4772 <= tmp_ivl_4774 & tmp_ivl_4769;
  tmp_ivl_4777 <= state_in_s1(153);
  tmp_ivl_4779 <= state_in_s0(153);
  tmp_ivl_4780 <= tmp_ivl_4777 & tmp_ivl_4779;
  LPM_q_ivl_4783 <= tmp_ivl_4785 & tmp_ivl_4780;
  new_AGEMA_signal_2753 <= tmp_ivl_4787(1);
  n3266 <= tmp_ivl_4787(0);
  tmp_ivl_4787 <= LPM_d0_ivl_4791(0 + 1 downto 0);
  tmp_ivl_4793 <= state_in_s1(169);
  tmp_ivl_4795 <= state_in_s0(169);
  tmp_ivl_4796 <= tmp_ivl_4793 & tmp_ivl_4795;
  LPM_q_ivl_4799 <= tmp_ivl_4801 & tmp_ivl_4796;
  tmp_ivl_4804 <= state_in_s1(105);
  tmp_ivl_4806 <= state_in_s0(105);
  tmp_ivl_4807 <= tmp_ivl_4804 & tmp_ivl_4806;
  LPM_q_ivl_4810 <= tmp_ivl_4812 & tmp_ivl_4807;
  new_AGEMA_signal_2755 <= tmp_ivl_4814(1);
  n3282 <= tmp_ivl_4814(0);
  tmp_ivl_4814 <= LPM_d0_ivl_4818(0 + 1 downto 0);
  tmp_ivl_4820 <= state_in_s1(90);
  tmp_ivl_4822 <= state_in_s0(90);
  tmp_ivl_4823 <= tmp_ivl_4820 & tmp_ivl_4822;
  LPM_q_ivl_4826 <= tmp_ivl_4828 & tmp_ivl_4823;
  tmp_ivl_4831 <= state_in_s1(154);
  tmp_ivl_4833 <= state_in_s0(154);
  tmp_ivl_4834 <= tmp_ivl_4831 & tmp_ivl_4833;
  LPM_q_ivl_4837 <= tmp_ivl_4839 & tmp_ivl_4834;
  new_AGEMA_signal_2758 <= tmp_ivl_4841(1);
  n3265 <= tmp_ivl_4841(0);
  tmp_ivl_4841 <= LPM_d0_ivl_4845(0 + 1 downto 0);
  tmp_ivl_4847 <= state_in_s1(106);
  tmp_ivl_4849 <= state_in_s0(106);
  tmp_ivl_4850 <= tmp_ivl_4847 & tmp_ivl_4849;
  LPM_q_ivl_4853 <= tmp_ivl_4855 & tmp_ivl_4850;
  tmp_ivl_4858 <= state_in_s1(170);
  tmp_ivl_4860 <= state_in_s0(170);
  tmp_ivl_4861 <= tmp_ivl_4858 & tmp_ivl_4860;
  LPM_q_ivl_4864 <= tmp_ivl_4866 & tmp_ivl_4861;
  new_AGEMA_signal_2760 <= tmp_ivl_4868(1);
  n3281 <= tmp_ivl_4868(0);
  tmp_ivl_4868 <= LPM_d0_ivl_4872(0 + 1 downto 0);
  tmp_ivl_4874 <= state_in_s1(91);
  tmp_ivl_4876 <= state_in_s0(91);
  tmp_ivl_4877 <= tmp_ivl_4874 & tmp_ivl_4876;
  LPM_q_ivl_4880 <= tmp_ivl_4882 & tmp_ivl_4877;
  tmp_ivl_4885 <= state_in_s1(155);
  tmp_ivl_4887 <= state_in_s0(155);
  tmp_ivl_4888 <= tmp_ivl_4885 & tmp_ivl_4887;
  LPM_q_ivl_4891 <= tmp_ivl_4893 & tmp_ivl_4888;
  new_AGEMA_signal_2763 <= tmp_ivl_4895(1);
  n3264 <= tmp_ivl_4895(0);
  tmp_ivl_4895 <= LPM_d0_ivl_4899(0 + 1 downto 0);
  tmp_ivl_4901 <= state_in_s1(92);
  tmp_ivl_4903 <= state_in_s0(92);
  tmp_ivl_4904 <= tmp_ivl_4901 & tmp_ivl_4903;
  LPM_q_ivl_4907 <= tmp_ivl_4909 & tmp_ivl_4904;
  tmp_ivl_4912 <= state_in_s1(156);
  tmp_ivl_4914 <= state_in_s0(156);
  tmp_ivl_4915 <= tmp_ivl_4912 & tmp_ivl_4914;
  LPM_q_ivl_4918 <= tmp_ivl_4920 & tmp_ivl_4915;
  new_AGEMA_signal_2766 <= tmp_ivl_4922(1);
  n3263 <= tmp_ivl_4922(0);
  tmp_ivl_4922 <= LPM_d0_ivl_4926(0 + 1 downto 0);
  tmp_ivl_4928 <= state_in_s1(93);
  tmp_ivl_4930 <= state_in_s0(93);
  tmp_ivl_4931 <= tmp_ivl_4928 & tmp_ivl_4930;
  LPM_q_ivl_4934 <= tmp_ivl_4936 & tmp_ivl_4931;
  tmp_ivl_4939 <= state_in_s1(157);
  tmp_ivl_4941 <= state_in_s0(157);
  tmp_ivl_4942 <= tmp_ivl_4939 & tmp_ivl_4941;
  LPM_q_ivl_4945 <= tmp_ivl_4947 & tmp_ivl_4942;
  new_AGEMA_signal_2769 <= tmp_ivl_4949(1);
  n3262 <= tmp_ivl_4949(0);
  tmp_ivl_4949 <= LPM_d0_ivl_4953(0 + 1 downto 0);
  tmp_ivl_4955 <= state_in_s1(94);
  tmp_ivl_4957 <= state_in_s0(94);
  tmp_ivl_4958 <= tmp_ivl_4955 & tmp_ivl_4957;
  LPM_q_ivl_4961 <= tmp_ivl_4963 & tmp_ivl_4958;
  tmp_ivl_4966 <= state_in_s1(158);
  tmp_ivl_4968 <= state_in_s0(158);
  tmp_ivl_4969 <= tmp_ivl_4966 & tmp_ivl_4968;
  LPM_q_ivl_4972 <= tmp_ivl_4974 & tmp_ivl_4969;
  new_AGEMA_signal_2772 <= tmp_ivl_4976(1);
  n3261 <= tmp_ivl_4976(0);
  tmp_ivl_4976 <= LPM_d0_ivl_4980(0 + 1 downto 0);
  tmp_ivl_4982 <= state_in_s1(95);
  tmp_ivl_4984 <= state_in_s0(95);
  tmp_ivl_4985 <= tmp_ivl_4982 & tmp_ivl_4984;
  LPM_q_ivl_4988 <= tmp_ivl_4990 & tmp_ivl_4985;
  tmp_ivl_4993 <= state_in_s1(159);
  tmp_ivl_4995 <= state_in_s0(159);
  tmp_ivl_4996 <= tmp_ivl_4993 & tmp_ivl_4995;
  LPM_q_ivl_4999 <= tmp_ivl_5001 & tmp_ivl_4996;
  new_AGEMA_signal_2775 <= tmp_ivl_5003(1);
  n3260 <= tmp_ivl_5003(0);
  tmp_ivl_5003 <= LPM_d0_ivl_5007(0 + 1 downto 0);
  tmp_ivl_5009 <= state_in_s1(80);
  tmp_ivl_5011 <= state_in_s0(80);
  tmp_ivl_5012 <= tmp_ivl_5009 & tmp_ivl_5011;
  LPM_q_ivl_5015 <= tmp_ivl_5017 & tmp_ivl_5012;
  tmp_ivl_5020 <= state_in_s1(144);
  tmp_ivl_5022 <= state_in_s0(144);
  tmp_ivl_5023 <= tmp_ivl_5020 & tmp_ivl_5022;
  LPM_q_ivl_5026 <= tmp_ivl_5028 & tmp_ivl_5023;
  new_AGEMA_signal_2778 <= tmp_ivl_5030(1);
  n3259 <= tmp_ivl_5030(0);
  tmp_ivl_5030 <= LPM_d0_ivl_5034(0 + 1 downto 0);
  tmp_ivl_5036 <= state_in_s1(81);
  tmp_ivl_5038 <= state_in_s0(81);
  tmp_ivl_5039 <= tmp_ivl_5036 & tmp_ivl_5038;
  LPM_q_ivl_5042 <= tmp_ivl_5044 & tmp_ivl_5039;
  tmp_ivl_5047 <= state_in_s1(145);
  tmp_ivl_5049 <= state_in_s0(145);
  tmp_ivl_5050 <= tmp_ivl_5047 & tmp_ivl_5049;
  LPM_q_ivl_5053 <= tmp_ivl_5055 & tmp_ivl_5050;
  new_AGEMA_signal_2780 <= tmp_ivl_5057(1);
  n3258 <= tmp_ivl_5057(0);
  tmp_ivl_5057 <= LPM_d0_ivl_5061(0 + 1 downto 0);
  tmp_ivl_5063 <= state_in_s1(82);
  tmp_ivl_5065 <= state_in_s0(82);
  tmp_ivl_5066 <= tmp_ivl_5063 & tmp_ivl_5065;
  LPM_q_ivl_5069 <= tmp_ivl_5071 & tmp_ivl_5066;
  tmp_ivl_5074 <= state_in_s1(146);
  tmp_ivl_5076 <= state_in_s0(146);
  tmp_ivl_5077 <= tmp_ivl_5074 & tmp_ivl_5076;
  LPM_q_ivl_5080 <= tmp_ivl_5082 & tmp_ivl_5077;
  new_AGEMA_signal_2783 <= tmp_ivl_5084(1);
  n3257 <= tmp_ivl_5084(0);
  tmp_ivl_5084 <= LPM_d0_ivl_5088(0 + 1 downto 0);
  tmp_ivl_5090 <= state_in_s1(83);
  tmp_ivl_5092 <= state_in_s0(83);
  tmp_ivl_5093 <= tmp_ivl_5090 & tmp_ivl_5092;
  LPM_q_ivl_5096 <= tmp_ivl_5098 & tmp_ivl_5093;
  tmp_ivl_5101 <= state_in_s1(147);
  tmp_ivl_5103 <= state_in_s0(147);
  tmp_ivl_5104 <= tmp_ivl_5101 & tmp_ivl_5103;
  LPM_q_ivl_5107 <= tmp_ivl_5109 & tmp_ivl_5104;
  new_AGEMA_signal_2786 <= tmp_ivl_5111(1);
  n3256 <= tmp_ivl_5111(0);
  tmp_ivl_5111 <= LPM_d0_ivl_5115(0 + 1 downto 0);
  tmp_ivl_5117 <= state_in_s1(84);
  tmp_ivl_5119 <= state_in_s0(84);
  tmp_ivl_5120 <= tmp_ivl_5117 & tmp_ivl_5119;
  LPM_q_ivl_5123 <= tmp_ivl_5125 & tmp_ivl_5120;
  tmp_ivl_5128 <= state_in_s1(148);
  tmp_ivl_5130 <= state_in_s0(148);
  tmp_ivl_5131 <= tmp_ivl_5128 & tmp_ivl_5130;
  LPM_q_ivl_5134 <= tmp_ivl_5136 & tmp_ivl_5131;
  new_AGEMA_signal_2788 <= tmp_ivl_5138(1);
  n3255 <= tmp_ivl_5138(0);
  tmp_ivl_5138 <= LPM_d0_ivl_5142(0 + 1 downto 0);
  tmp_ivl_5144 <= state_in_s1(85);
  tmp_ivl_5146 <= state_in_s0(85);
  tmp_ivl_5147 <= tmp_ivl_5144 & tmp_ivl_5146;
  LPM_q_ivl_5150 <= tmp_ivl_5152 & tmp_ivl_5147;
  tmp_ivl_5155 <= state_in_s1(149);
  tmp_ivl_5157 <= state_in_s0(149);
  tmp_ivl_5158 <= tmp_ivl_5155 & tmp_ivl_5157;
  LPM_q_ivl_5161 <= tmp_ivl_5163 & tmp_ivl_5158;
  new_AGEMA_signal_2790 <= tmp_ivl_5165(1);
  n3254 <= tmp_ivl_5165(0);
  tmp_ivl_5165 <= LPM_d0_ivl_5169(0 + 1 downto 0);
  tmp_ivl_5171 <= state_in_s1(86);
  tmp_ivl_5173 <= state_in_s0(86);
  tmp_ivl_5174 <= tmp_ivl_5171 & tmp_ivl_5173;
  LPM_q_ivl_5177 <= tmp_ivl_5179 & tmp_ivl_5174;
  tmp_ivl_5182 <= state_in_s1(150);
  tmp_ivl_5184 <= state_in_s0(150);
  tmp_ivl_5185 <= tmp_ivl_5182 & tmp_ivl_5184;
  LPM_q_ivl_5188 <= tmp_ivl_5190 & tmp_ivl_5185;
  new_AGEMA_signal_2793 <= tmp_ivl_5192(1);
  n3253 <= tmp_ivl_5192(0);
  tmp_ivl_5192 <= LPM_d0_ivl_5196(0 + 1 downto 0);
  tmp_ivl_5198 <= state_in_s1(87);
  tmp_ivl_5200 <= state_in_s0(87);
  tmp_ivl_5201 <= tmp_ivl_5198 & tmp_ivl_5200;
  LPM_q_ivl_5204 <= tmp_ivl_5206 & tmp_ivl_5201;
  tmp_ivl_5209 <= state_in_s1(151);
  tmp_ivl_5211 <= state_in_s0(151);
  tmp_ivl_5212 <= tmp_ivl_5209 & tmp_ivl_5211;
  LPM_q_ivl_5215 <= tmp_ivl_5217 & tmp_ivl_5212;
  new_AGEMA_signal_2795 <= tmp_ivl_5219(1);
  n3252 <= tmp_ivl_5219(0);
  tmp_ivl_5219 <= LPM_d0_ivl_5223(0 + 1 downto 0);
  tmp_ivl_5225 <= state_in_s1(72);
  tmp_ivl_5227 <= state_in_s0(72);
  tmp_ivl_5228 <= tmp_ivl_5225 & tmp_ivl_5227;
  LPM_q_ivl_5231 <= tmp_ivl_5233 & tmp_ivl_5228;
  tmp_ivl_5236 <= state_in_s1(136);
  tmp_ivl_5238 <= state_in_s0(136);
  tmp_ivl_5239 <= tmp_ivl_5236 & tmp_ivl_5238;
  LPM_q_ivl_5242 <= tmp_ivl_5244 & tmp_ivl_5239;
  new_AGEMA_signal_2797 <= tmp_ivl_5246(1);
  n3251 <= tmp_ivl_5246(0);
  tmp_ivl_5246 <= LPM_d0_ivl_5250(0 + 1 downto 0);
  tmp_ivl_5252 <= state_in_s1(137);
  tmp_ivl_5254 <= state_in_s0(137);
  tmp_ivl_5255 <= tmp_ivl_5252 & tmp_ivl_5254;
  LPM_q_ivl_5258 <= tmp_ivl_5260 & tmp_ivl_5255;
  tmp_ivl_5263 <= state_in_s1(73);
  tmp_ivl_5265 <= state_in_s0(73);
  tmp_ivl_5266 <= tmp_ivl_5263 & tmp_ivl_5265;
  LPM_q_ivl_5269 <= tmp_ivl_5271 & tmp_ivl_5266;
  new_AGEMA_signal_2800 <= tmp_ivl_5273(1);
  n3250 <= tmp_ivl_5273(0);
  tmp_ivl_5273 <= LPM_d0_ivl_5277(0 + 1 downto 0);
  tmp_ivl_5279 <= state_in_s1(138);
  tmp_ivl_5281 <= state_in_s0(138);
  tmp_ivl_5282 <= tmp_ivl_5279 & tmp_ivl_5281;
  LPM_q_ivl_5285 <= tmp_ivl_5287 & tmp_ivl_5282;
  tmp_ivl_5290 <= state_in_s1(74);
  tmp_ivl_5292 <= state_in_s0(74);
  tmp_ivl_5293 <= tmp_ivl_5290 & tmp_ivl_5292;
  LPM_q_ivl_5296 <= tmp_ivl_5298 & tmp_ivl_5293;
  new_AGEMA_signal_2803 <= tmp_ivl_5300(1);
  n3249 <= tmp_ivl_5300(0);
  tmp_ivl_5300 <= LPM_d0_ivl_5304(0 + 1 downto 0);
  tmp_ivl_5306 <= state_in_s1(75);
  tmp_ivl_5308 <= state_in_s0(75);
  tmp_ivl_5309 <= tmp_ivl_5306 & tmp_ivl_5308;
  LPM_q_ivl_5312 <= tmp_ivl_5314 & tmp_ivl_5309;
  tmp_ivl_5317 <= state_in_s1(139);
  tmp_ivl_5319 <= state_in_s0(139);
  tmp_ivl_5320 <= tmp_ivl_5317 & tmp_ivl_5319;
  LPM_q_ivl_5323 <= tmp_ivl_5325 & tmp_ivl_5320;
  new_AGEMA_signal_2805 <= tmp_ivl_5327(1);
  n3248 <= tmp_ivl_5327(0);
  tmp_ivl_5327 <= LPM_d0_ivl_5331(0 + 1 downto 0);
  tmp_ivl_5333 <= state_in_s1(76);
  tmp_ivl_5335 <= state_in_s0(76);
  tmp_ivl_5336 <= tmp_ivl_5333 & tmp_ivl_5335;
  LPM_q_ivl_5339 <= tmp_ivl_5341 & tmp_ivl_5336;
  tmp_ivl_5344 <= state_in_s1(140);
  tmp_ivl_5346 <= state_in_s0(140);
  tmp_ivl_5347 <= tmp_ivl_5344 & tmp_ivl_5346;
  LPM_q_ivl_5350 <= tmp_ivl_5352 & tmp_ivl_5347;
  new_AGEMA_signal_2807 <= tmp_ivl_5354(1);
  n3247 <= tmp_ivl_5354(0);
  tmp_ivl_5354 <= LPM_d0_ivl_5358(0 + 1 downto 0);
  tmp_ivl_5360 <= state_in_s1(141);
  tmp_ivl_5362 <= state_in_s0(141);
  tmp_ivl_5363 <= tmp_ivl_5360 & tmp_ivl_5362;
  LPM_q_ivl_5366 <= tmp_ivl_5368 & tmp_ivl_5363;
  tmp_ivl_5371 <= state_in_s1(77);
  tmp_ivl_5373 <= state_in_s0(77);
  tmp_ivl_5374 <= tmp_ivl_5371 & tmp_ivl_5373;
  LPM_q_ivl_5377 <= tmp_ivl_5379 & tmp_ivl_5374;
  new_AGEMA_signal_2810 <= tmp_ivl_5381(1);
  n3246 <= tmp_ivl_5381(0);
  tmp_ivl_5381 <= LPM_d0_ivl_5385(0 + 1 downto 0);
  tmp_ivl_5387 <= state_in_s1(142);
  tmp_ivl_5389 <= state_in_s0(142);
  tmp_ivl_5390 <= tmp_ivl_5387 & tmp_ivl_5389;
  LPM_q_ivl_5393 <= tmp_ivl_5395 & tmp_ivl_5390;
  tmp_ivl_5398 <= state_in_s1(78);
  tmp_ivl_5400 <= state_in_s0(78);
  tmp_ivl_5401 <= tmp_ivl_5398 & tmp_ivl_5400;
  LPM_q_ivl_5404 <= tmp_ivl_5406 & tmp_ivl_5401;
  new_AGEMA_signal_2813 <= tmp_ivl_5408(1);
  n3245 <= tmp_ivl_5408(0);
  tmp_ivl_5408 <= LPM_d0_ivl_5412(0 + 1 downto 0);
  tmp_ivl_5414 <= state_in_s1(79);
  tmp_ivl_5416 <= state_in_s0(79);
  tmp_ivl_5417 <= tmp_ivl_5414 & tmp_ivl_5416;
  LPM_q_ivl_5420 <= tmp_ivl_5422 & tmp_ivl_5417;
  tmp_ivl_5425 <= state_in_s1(143);
  tmp_ivl_5427 <= state_in_s0(143);
  tmp_ivl_5428 <= tmp_ivl_5425 & tmp_ivl_5427;
  LPM_q_ivl_5431 <= tmp_ivl_5433 & tmp_ivl_5428;
  new_AGEMA_signal_2816 <= tmp_ivl_5435(1);
  n3244 <= tmp_ivl_5435(0);
  tmp_ivl_5435 <= LPM_d0_ivl_5439(0 + 1 downto 0);
  tmp_ivl_5441 <= state_in_s1(128);
  tmp_ivl_5443 <= state_in_s0(128);
  tmp_ivl_5444 <= tmp_ivl_5441 & tmp_ivl_5443;
  LPM_q_ivl_5447 <= tmp_ivl_5449 & tmp_ivl_5444;
  tmp_ivl_5452 <= state_in_s1(64);
  tmp_ivl_5454 <= state_in_s0(64);
  tmp_ivl_5455 <= tmp_ivl_5452 & tmp_ivl_5454;
  LPM_q_ivl_5458 <= tmp_ivl_5460 & tmp_ivl_5455;
  new_AGEMA_signal_2819 <= tmp_ivl_5462(1);
  n3243 <= tmp_ivl_5462(0);
  tmp_ivl_5462 <= LPM_d0_ivl_5466(0 + 1 downto 0);
  tmp_ivl_5468 <= state_in_s1(129);
  tmp_ivl_5470 <= state_in_s0(129);
  tmp_ivl_5471 <= tmp_ivl_5468 & tmp_ivl_5470;
  LPM_q_ivl_5474 <= tmp_ivl_5476 & tmp_ivl_5471;
  tmp_ivl_5479 <= state_in_s1(65);
  tmp_ivl_5481 <= state_in_s0(65);
  tmp_ivl_5482 <= tmp_ivl_5479 & tmp_ivl_5481;
  LPM_q_ivl_5485 <= tmp_ivl_5487 & tmp_ivl_5482;
  new_AGEMA_signal_2821 <= tmp_ivl_5489(1);
  n3242 <= tmp_ivl_5489(0);
  tmp_ivl_5489 <= LPM_d0_ivl_5493(0 + 1 downto 0);
  tmp_ivl_5495 <= state_in_s1(66);
  tmp_ivl_5497 <= state_in_s0(66);
  tmp_ivl_5498 <= tmp_ivl_5495 & tmp_ivl_5497;
  LPM_q_ivl_5501 <= tmp_ivl_5503 & tmp_ivl_5498;
  tmp_ivl_5506 <= state_in_s1(130);
  tmp_ivl_5508 <= state_in_s0(130);
  tmp_ivl_5509 <= tmp_ivl_5506 & tmp_ivl_5508;
  LPM_q_ivl_5512 <= tmp_ivl_5514 & tmp_ivl_5509;
  new_AGEMA_signal_2823 <= tmp_ivl_5516(1);
  n3241 <= tmp_ivl_5516(0);
  tmp_ivl_5516 <= LPM_d0_ivl_5520(0 + 1 downto 0);
  tmp_ivl_5522 <= state_in_s1(131);
  tmp_ivl_5524 <= state_in_s0(131);
  tmp_ivl_5525 <= tmp_ivl_5522 & tmp_ivl_5524;
  LPM_q_ivl_5528 <= tmp_ivl_5530 & tmp_ivl_5525;
  tmp_ivl_5533 <= state_in_s1(67);
  tmp_ivl_5535 <= state_in_s0(67);
  tmp_ivl_5536 <= tmp_ivl_5533 & tmp_ivl_5535;
  LPM_q_ivl_5539 <= tmp_ivl_5541 & tmp_ivl_5536;
  new_AGEMA_signal_2825 <= tmp_ivl_5543(1);
  n3240 <= tmp_ivl_5543(0);
  tmp_ivl_5543 <= LPM_d0_ivl_5547(0 + 1 downto 0);
  tmp_ivl_5549 <= state_in_s1(132);
  tmp_ivl_5551 <= state_in_s0(132);
  tmp_ivl_5552 <= tmp_ivl_5549 & tmp_ivl_5551;
  LPM_q_ivl_5555 <= tmp_ivl_5557 & tmp_ivl_5552;
  tmp_ivl_5560 <= state_in_s1(68);
  tmp_ivl_5562 <= state_in_s0(68);
  tmp_ivl_5563 <= tmp_ivl_5560 & tmp_ivl_5562;
  LPM_q_ivl_5566 <= tmp_ivl_5568 & tmp_ivl_5563;
  new_AGEMA_signal_2828 <= tmp_ivl_5570(1);
  n3238 <= tmp_ivl_5570(0);
  tmp_ivl_5570 <= LPM_d0_ivl_5574(0 + 1 downto 0);
  tmp_ivl_5576 <= state_in_s1(184);
  tmp_ivl_5578 <= state_in_s0(184);
  tmp_ivl_5579 <= tmp_ivl_5576 & tmp_ivl_5578;
  LPM_q_ivl_5582 <= tmp_ivl_5584 & tmp_ivl_5579;
  tmp_ivl_5587 <= state_in_s1(120);
  tmp_ivl_5589 <= state_in_s0(120);
  tmp_ivl_5590 <= tmp_ivl_5587 & tmp_ivl_5589;
  LPM_q_ivl_5593 <= tmp_ivl_5595 & tmp_ivl_5590;
  new_AGEMA_signal_2831 <= tmp_ivl_5597(1);
  n4041 <= tmp_ivl_5597(0);
  tmp_ivl_5597 <= LPM_d0_ivl_5601(0 + 1 downto 0);
  LPM_q_ivl_5602 <= rcon(0);
  tmp_ivl_5604 <= new_AGEMA_signal_2831 & n4041;
  LPM_q_ivl_5607 <= tmp_ivl_5609 & tmp_ivl_5604;
  tmp_ivl_5613 <= tmp_ivl_5611 & n4068;
  LPM_q_ivl_5616 <= tmp_ivl_5618 & tmp_ivl_5613;
  new_AGEMA_signal_2989 <= tmp_ivl_5622(1);
  tmp_ivl_5620 <= tmp_ivl_5622(0);
  tmp_ivl_5622 <= LPM_d0_ivl_5626(0 + 1 downto 0);
  tmp_ivl_5628 <= state_in_s1(176);
  tmp_ivl_5630 <= state_in_s0(176);
  tmp_ivl_5631 <= tmp_ivl_5628 & tmp_ivl_5630;
  LPM_q_ivl_5634 <= tmp_ivl_5636 & tmp_ivl_5631;
  tmp_ivl_5639 <= state_in_s1(112);
  tmp_ivl_5641 <= state_in_s0(112);
  tmp_ivl_5642 <= tmp_ivl_5639 & tmp_ivl_5641;
  LPM_q_ivl_5645 <= tmp_ivl_5647 & tmp_ivl_5642;
  new_AGEMA_signal_2834 <= tmp_ivl_5649(1);
  n3237 <= tmp_ivl_5649(0);
  tmp_ivl_5649 <= LPM_d0_ivl_5653(0 + 1 downto 0);
  tmp_ivl_5655 <= state_in_s1(133);
  tmp_ivl_5657 <= state_in_s0(133);
  tmp_ivl_5658 <= tmp_ivl_5655 & tmp_ivl_5657;
  LPM_q_ivl_5661 <= tmp_ivl_5663 & tmp_ivl_5658;
  tmp_ivl_5666 <= state_in_s1(69);
  tmp_ivl_5668 <= state_in_s0(69);
  tmp_ivl_5669 <= tmp_ivl_5666 & tmp_ivl_5668;
  LPM_q_ivl_5672 <= tmp_ivl_5674 & tmp_ivl_5669;
  new_AGEMA_signal_2837 <= tmp_ivl_5676(1);
  n3236 <= tmp_ivl_5676(0);
  tmp_ivl_5676 <= LPM_d0_ivl_5680(0 + 1 downto 0);
  tmp_ivl_5682 <= state_in_s1(134);
  tmp_ivl_5684 <= state_in_s0(134);
  tmp_ivl_5685 <= tmp_ivl_5682 & tmp_ivl_5684;
  LPM_q_ivl_5688 <= tmp_ivl_5690 & tmp_ivl_5685;
  tmp_ivl_5693 <= state_in_s1(70);
  tmp_ivl_5695 <= state_in_s0(70);
  tmp_ivl_5696 <= tmp_ivl_5693 & tmp_ivl_5695;
  LPM_q_ivl_5699 <= tmp_ivl_5701 & tmp_ivl_5696;
  new_AGEMA_signal_2840 <= tmp_ivl_5703(1);
  n3235 <= tmp_ivl_5703(0);
  tmp_ivl_5703 <= LPM_d0_ivl_5707(0 + 1 downto 0);
  tmp_ivl_5709 <= state_in_s1(188);
  tmp_ivl_5711 <= state_in_s0(188);
  tmp_ivl_5712 <= tmp_ivl_5709 & tmp_ivl_5711;
  LPM_q_ivl_5715 <= tmp_ivl_5717 & tmp_ivl_5712;
  tmp_ivl_5720 <= state_in_s1(124);
  tmp_ivl_5722 <= state_in_s0(124);
  tmp_ivl_5723 <= tmp_ivl_5720 & tmp_ivl_5722;
  LPM_q_ivl_5726 <= tmp_ivl_5728 & tmp_ivl_5723;
  new_AGEMA_signal_2843 <= tmp_ivl_5730(1);
  n4208 <= tmp_ivl_5730(0);
  tmp_ivl_5730 <= LPM_d0_ivl_5734(0 + 1 downto 0);
  tmp_ivl_5738 <= rcon(0);
  tmp_ivl_5739 <= tmp_ivl_5735 & tmp_ivl_5738;
  LPM_q_ivl_5742 <= tmp_ivl_5744 & tmp_ivl_5739;
  tmp_ivl_5746 <= new_AGEMA_signal_2843 & n4208;
  LPM_q_ivl_5749 <= tmp_ivl_5751 & tmp_ivl_5746;
  new_AGEMA_signal_2990 <= tmp_ivl_5753(1);
  n3232 <= tmp_ivl_5753(0);
  tmp_ivl_5753 <= LPM_d0_ivl_5757(0 + 1 downto 0);
  tmp_ivl_5759 <= state_in_s1(135);
  tmp_ivl_5761 <= state_in_s0(135);
  tmp_ivl_5762 <= tmp_ivl_5759 & tmp_ivl_5761;
  LPM_q_ivl_5765 <= tmp_ivl_5767 & tmp_ivl_5762;
  tmp_ivl_5770 <= state_in_s1(71);
  tmp_ivl_5772 <= state_in_s0(71);
  tmp_ivl_5773 <= tmp_ivl_5770 & tmp_ivl_5772;
  LPM_q_ivl_5776 <= tmp_ivl_5778 & tmp_ivl_5773;
  new_AGEMA_signal_2846 <= tmp_ivl_5780(1);
  n3234 <= tmp_ivl_5780(0);
  tmp_ivl_5780 <= LPM_d0_ivl_5784(0 + 1 downto 0);
  LPM_q_ivl_5785 <= rcon(1);
  LPM_q_ivl_5787 <= rcon(0);
  tmp_ivl_5790 <= state_in_s1(185);
  tmp_ivl_5792 <= state_in_s0(185);
  tmp_ivl_5793 <= tmp_ivl_5790 & tmp_ivl_5792;
  LPM_q_ivl_5796 <= tmp_ivl_5798 & tmp_ivl_5793;
  tmp_ivl_5801 <= state_in_s1(121);
  tmp_ivl_5803 <= state_in_s0(121);
  tmp_ivl_5804 <= tmp_ivl_5801 & tmp_ivl_5803;
  LPM_q_ivl_5807 <= tmp_ivl_5809 & tmp_ivl_5804;
  new_AGEMA_signal_2849 <= tmp_ivl_5811(1);
  n4066 <= tmp_ivl_5811(0);
  tmp_ivl_5811 <= LPM_d0_ivl_5815(0 + 1 downto 0);
  tmp_ivl_5818 <= tmp_ivl_5816 & n4206;
  LPM_q_ivl_5821 <= tmp_ivl_5823 & tmp_ivl_5818;
  tmp_ivl_5825 <= new_AGEMA_signal_2849 & n4066;
  LPM_q_ivl_5828 <= tmp_ivl_5830 & tmp_ivl_5825;
  new_AGEMA_signal_3513 <= tmp_ivl_5834(1);
  tmp_ivl_5832 <= tmp_ivl_5834(0);
  tmp_ivl_5834 <= LPM_d0_ivl_5838(0 + 1 downto 0);
  tmp_ivl_5840 <= state_in_s1(186);
  tmp_ivl_5842 <= state_in_s0(186);
  tmp_ivl_5843 <= tmp_ivl_5840 & tmp_ivl_5842;
  LPM_q_ivl_5846 <= tmp_ivl_5848 & tmp_ivl_5843;
  tmp_ivl_5851 <= state_in_s1(122);
  tmp_ivl_5853 <= state_in_s0(122);
  tmp_ivl_5854 <= tmp_ivl_5851 & tmp_ivl_5853;
  LPM_q_ivl_5857 <= tmp_ivl_5859 & tmp_ivl_5854;
  new_AGEMA_signal_2852 <= tmp_ivl_5861(1);
  n4069 <= tmp_ivl_5861(0);
  tmp_ivl_5861 <= LPM_d0_ivl_5865(0 + 1 downto 0);
  LPM_q_ivl_5866 <= rcon(2);
  tmp_ivl_5868 <= new_AGEMA_signal_2852 & n4069;
  LPM_q_ivl_5871 <= tmp_ivl_5873 & tmp_ivl_5868;
  tmp_ivl_5877 <= tmp_ivl_5875 & n4087;
  LPM_q_ivl_5880 <= tmp_ivl_5882 & tmp_ivl_5877;
  new_AGEMA_signal_3824 <= tmp_ivl_5884(1);
  n3287 <= tmp_ivl_5884(0);
  tmp_ivl_5884 <= LPM_d0_ivl_5888(0 + 1 downto 0);
  LPM_q_ivl_5889 <= rcon(2);
  LPM_q_ivl_5891 <= rcon(3);
  tmp_ivl_5895 <= tmp_ivl_5893 & n4084;
  LPM_q_ivl_5898 <= tmp_ivl_5900 & tmp_ivl_5895;
  tmp_ivl_5903 <= state_in_s1(187);
  tmp_ivl_5905 <= state_in_s0(187);
  tmp_ivl_5906 <= tmp_ivl_5903 & tmp_ivl_5905;
  LPM_q_ivl_5909 <= tmp_ivl_5911 & tmp_ivl_5906;
  new_AGEMA_signal_4140 <= tmp_ivl_5913(1);
  n4081 <= tmp_ivl_5913(0);
  tmp_ivl_5913 <= LPM_d0_ivl_5917(0 + 1 downto 0);
  tmp_ivl_5919 <= state_in_s1(123);
  tmp_ivl_5921 <= state_in_s0(123);
  tmp_ivl_5922 <= tmp_ivl_5919 & tmp_ivl_5921;
  LPM_q_ivl_5925 <= tmp_ivl_5927 & tmp_ivl_5922;
  tmp_ivl_5929 <= new_AGEMA_signal_4140 & n4081;
  LPM_q_ivl_5932 <= tmp_ivl_5934 & tmp_ivl_5929;
  new_AGEMA_signal_4432 <= tmp_ivl_5936(1);
  n3233 <= tmp_ivl_5936(0);
  tmp_ivl_5936 <= LPM_d0_ivl_5940(0 + 1 downto 0);
  tmp_ivl_5943 <= tmp_ivl_5941 & n4084;
  LPM_q_ivl_5946 <= tmp_ivl_5948 & tmp_ivl_5943;
  tmp_ivl_5951 <= state_in_s1(191);
  tmp_ivl_5953 <= state_in_s0(191);
  tmp_ivl_5954 <= tmp_ivl_5951 & tmp_ivl_5953;
  LPM_q_ivl_5957 <= tmp_ivl_5959 & tmp_ivl_5954;
  new_AGEMA_signal_4142 <= tmp_ivl_5961(1);
  n4085 <= tmp_ivl_5961(0);
  tmp_ivl_5961 <= LPM_d0_ivl_5965(0 + 1 downto 0);
  tmp_ivl_5966 <= new_AGEMA_signal_4142 & n4085;
  LPM_q_ivl_5969 <= tmp_ivl_5971 & tmp_ivl_5966;
  tmp_ivl_5974 <= state_in_s1(127);
  tmp_ivl_5976 <= state_in_s0(127);
  tmp_ivl_5977 <= tmp_ivl_5974 & tmp_ivl_5976;
  LPM_q_ivl_5980 <= tmp_ivl_5982 & tmp_ivl_5977;
  new_AGEMA_signal_4433 <= tmp_ivl_5984(1);
  n3239 <= tmp_ivl_5984(0);
  tmp_ivl_5984 <= LPM_d0_ivl_5988(0 + 1 downto 0);
  tmp_ivl_5990 <= state_in_s1(190);
  tmp_ivl_5992 <= state_in_s0(190);
  tmp_ivl_5993 <= tmp_ivl_5990 & tmp_ivl_5992;
  LPM_q_ivl_5996 <= tmp_ivl_5998 & tmp_ivl_5993;
  tmp_ivl_6001 <= state_in_s1(126);
  tmp_ivl_6003 <= state_in_s0(126);
  tmp_ivl_6004 <= tmp_ivl_6001 & tmp_ivl_6003;
  LPM_q_ivl_6007 <= tmp_ivl_6009 & tmp_ivl_6004;
  new_AGEMA_signal_2855 <= tmp_ivl_6011(1);
  n4086 <= tmp_ivl_6011(0);
  tmp_ivl_6011 <= LPM_d0_ivl_6015(0 + 1 downto 0);
  tmp_ivl_6018 <= tmp_ivl_6016 & n4087;
  LPM_q_ivl_6021 <= tmp_ivl_6023 & tmp_ivl_6018;
  tmp_ivl_6025 <= new_AGEMA_signal_2855 & n4086;
  LPM_q_ivl_6028 <= tmp_ivl_6030 & tmp_ivl_6025;
  new_AGEMA_signal_3826 <= tmp_ivl_6032(1);
  n3230 <= tmp_ivl_6032(0);
  tmp_ivl_6032 <= LPM_d0_ivl_6036(0 + 1 downto 0);
  tmp_ivl_6038 <= state_in_s1(125);
  tmp_ivl_6040 <= state_in_s0(125);
  tmp_ivl_6041 <= tmp_ivl_6038 & tmp_ivl_6040;
  LPM_q_ivl_6044 <= tmp_ivl_6046 & tmp_ivl_6041;
  tmp_ivl_6049 <= state_in_s1(189);
  tmp_ivl_6051 <= state_in_s0(189);
  tmp_ivl_6052 <= tmp_ivl_6049 & tmp_ivl_6051;
  LPM_q_ivl_6055 <= tmp_ivl_6057 & tmp_ivl_6052;
  new_AGEMA_signal_2858 <= tmp_ivl_6059(1);
  n4103 <= tmp_ivl_6059(0);
  tmp_ivl_6059 <= LPM_d0_ivl_6063(0 + 1 downto 0);
  tmp_ivl_6066 <= tmp_ivl_6064 & n4206;
  LPM_q_ivl_6069 <= tmp_ivl_6071 & tmp_ivl_6066;
  tmp_ivl_6073 <= new_AGEMA_signal_2858 & n4103;
  LPM_q_ivl_6076 <= tmp_ivl_6078 & tmp_ivl_6073;
  new_AGEMA_signal_3515 <= tmp_ivl_6080(1);
  n3231 <= tmp_ivl_6080(0);
  tmp_ivl_6080 <= LPM_d0_ivl_6084(0 + 1 downto 0);
  tmp_ivl_6086 <= y0(0);
  LPM_q_ivl_6088 <= new_AGEMA_signal_2655 & tmp_ivl_6086;
  new_AGEMA_signal_3047 <= LPM_d0_ivl_6090(1);
  SboxInst_n320 <= LPM_d0_ivl_6090(0);
  tmp_ivl_6093 <= y0(10);
  LPM_q_ivl_6095 <= new_AGEMA_signal_2653 & tmp_ivl_6093;
  new_AGEMA_signal_3048 <= LPM_d0_ivl_6097(1);
  SboxInst_n319 <= LPM_d0_ivl_6097(0);
  tmp_ivl_6100 <= y0(11);
  LPM_q_ivl_6102 <= new_AGEMA_signal_2651 & tmp_ivl_6100;
  new_AGEMA_signal_3049 <= LPM_d0_ivl_6104(1);
  SboxInst_n318 <= LPM_d0_ivl_6104(0);
  tmp_ivl_6107 <= y0(12);
  LPM_q_ivl_6109 <= new_AGEMA_signal_2649 & tmp_ivl_6107;
  new_AGEMA_signal_3050 <= LPM_d0_ivl_6111(1);
  SboxInst_n317 <= LPM_d0_ivl_6111(0);
  tmp_ivl_6114 <= y0(13);
  LPM_q_ivl_6116 <= new_AGEMA_signal_2647 & tmp_ivl_6114;
  new_AGEMA_signal_3051 <= LPM_d0_ivl_6118(1);
  SboxInst_n316 <= LPM_d0_ivl_6118(0);
  tmp_ivl_6121 <= y0(14);
  LPM_q_ivl_6123 <= new_AGEMA_signal_2645 & tmp_ivl_6121;
  new_AGEMA_signal_3052 <= LPM_d0_ivl_6125(1);
  SboxInst_n315 <= LPM_d0_ivl_6125(0);
  tmp_ivl_6128 <= y0(15);
  LPM_q_ivl_6130 <= new_AGEMA_signal_2643 & tmp_ivl_6128;
  new_AGEMA_signal_3053 <= LPM_d0_ivl_6132(1);
  SboxInst_n314 <= LPM_d0_ivl_6132(0);
  tmp_ivl_6135 <= y0(16);
  LPM_q_ivl_6137 <= new_AGEMA_signal_2641 & tmp_ivl_6135;
  new_AGEMA_signal_3054 <= LPM_d0_ivl_6139(1);
  SboxInst_n313 <= LPM_d0_ivl_6139(0);
  tmp_ivl_6142 <= y0(17);
  LPM_q_ivl_6144 <= new_AGEMA_signal_2639 & tmp_ivl_6142;
  new_AGEMA_signal_3055 <= LPM_d0_ivl_6146(1);
  SboxInst_n312 <= LPM_d0_ivl_6146(0);
  tmp_ivl_6149 <= y0(18);
  LPM_q_ivl_6151 <= new_AGEMA_signal_2637 & tmp_ivl_6149;
  new_AGEMA_signal_3056 <= LPM_d0_ivl_6153(1);
  SboxInst_n311 <= LPM_d0_ivl_6153(0);
  tmp_ivl_6156 <= y0(19);
  LPM_q_ivl_6158 <= new_AGEMA_signal_2635 & tmp_ivl_6156;
  new_AGEMA_signal_3057 <= LPM_d0_ivl_6160(1);
  SboxInst_n310 <= LPM_d0_ivl_6160(0);
  tmp_ivl_6163 <= y0(1);
  LPM_q_ivl_6165 <= new_AGEMA_signal_2633 & tmp_ivl_6163;
  new_AGEMA_signal_3058 <= LPM_d0_ivl_6167(1);
  SboxInst_n309 <= LPM_d0_ivl_6167(0);
  tmp_ivl_6170 <= y0(20);
  LPM_q_ivl_6172 <= new_AGEMA_signal_2631 & tmp_ivl_6170;
  new_AGEMA_signal_3059 <= LPM_d0_ivl_6174(1);
  SboxInst_n308 <= LPM_d0_ivl_6174(0);
  tmp_ivl_6177 <= y0(21);
  LPM_q_ivl_6179 <= new_AGEMA_signal_2629 & tmp_ivl_6177;
  new_AGEMA_signal_3060 <= LPM_d0_ivl_6181(1);
  SboxInst_n307 <= LPM_d0_ivl_6181(0);
  tmp_ivl_6184 <= y0(22);
  LPM_q_ivl_6186 <= new_AGEMA_signal_2627 & tmp_ivl_6184;
  new_AGEMA_signal_3061 <= LPM_d0_ivl_6188(1);
  SboxInst_n306 <= LPM_d0_ivl_6188(0);
  tmp_ivl_6191 <= y0(23);
  LPM_q_ivl_6193 <= new_AGEMA_signal_2625 & tmp_ivl_6191;
  new_AGEMA_signal_3062 <= LPM_d0_ivl_6195(1);
  SboxInst_n305 <= LPM_d0_ivl_6195(0);
  tmp_ivl_6198 <= y0(24);
  LPM_q_ivl_6200 <= new_AGEMA_signal_2623 & tmp_ivl_6198;
  new_AGEMA_signal_3063 <= LPM_d0_ivl_6202(1);
  SboxInst_n304 <= LPM_d0_ivl_6202(0);
  tmp_ivl_6205 <= y0(25);
  LPM_q_ivl_6207 <= new_AGEMA_signal_2621 & tmp_ivl_6205;
  new_AGEMA_signal_3064 <= LPM_d0_ivl_6209(1);
  SboxInst_n303 <= LPM_d0_ivl_6209(0);
  tmp_ivl_6212 <= y0(26);
  LPM_q_ivl_6214 <= new_AGEMA_signal_2619 & tmp_ivl_6212;
  new_AGEMA_signal_3065 <= LPM_d0_ivl_6216(1);
  SboxInst_n302 <= LPM_d0_ivl_6216(0);
  tmp_ivl_6219 <= y0(27);
  LPM_q_ivl_6221 <= new_AGEMA_signal_2617 & tmp_ivl_6219;
  new_AGEMA_signal_3066 <= LPM_d0_ivl_6223(1);
  SboxInst_n301 <= LPM_d0_ivl_6223(0);
  tmp_ivl_6226 <= y0(28);
  LPM_q_ivl_6228 <= new_AGEMA_signal_2615 & tmp_ivl_6226;
  new_AGEMA_signal_3067 <= LPM_d0_ivl_6230(1);
  SboxInst_n300 <= LPM_d0_ivl_6230(0);
  tmp_ivl_6233 <= y0(29);
  LPM_q_ivl_6235 <= new_AGEMA_signal_2613 & tmp_ivl_6233;
  new_AGEMA_signal_3068 <= LPM_d0_ivl_6237(1);
  SboxInst_n299 <= LPM_d0_ivl_6237(0);
  tmp_ivl_6240 <= y0(2);
  LPM_q_ivl_6242 <= new_AGEMA_signal_2611 & tmp_ivl_6240;
  new_AGEMA_signal_3069 <= LPM_d0_ivl_6244(1);
  SboxInst_n298 <= LPM_d0_ivl_6244(0);
  tmp_ivl_6247 <= y0(30);
  LPM_q_ivl_6249 <= new_AGEMA_signal_2609 & tmp_ivl_6247;
  new_AGEMA_signal_3070 <= LPM_d0_ivl_6251(1);
  SboxInst_n297 <= LPM_d0_ivl_6251(0);
  tmp_ivl_6254 <= y0(31);
  LPM_q_ivl_6256 <= new_AGEMA_signal_2607 & tmp_ivl_6254;
  new_AGEMA_signal_3071 <= LPM_d0_ivl_6258(1);
  SboxInst_n296 <= LPM_d0_ivl_6258(0);
  tmp_ivl_6261 <= y0(32);
  LPM_q_ivl_6263 <= new_AGEMA_signal_2605 & tmp_ivl_6261;
  new_AGEMA_signal_3072 <= LPM_d0_ivl_6265(1);
  SboxInst_n295 <= LPM_d0_ivl_6265(0);
  tmp_ivl_6268 <= y0(33);
  LPM_q_ivl_6270 <= new_AGEMA_signal_2603 & tmp_ivl_6268;
  new_AGEMA_signal_3073 <= LPM_d0_ivl_6272(1);
  SboxInst_n294 <= LPM_d0_ivl_6272(0);
  tmp_ivl_6275 <= y0(34);
  LPM_q_ivl_6277 <= new_AGEMA_signal_2601 & tmp_ivl_6275;
  new_AGEMA_signal_3074 <= LPM_d0_ivl_6279(1);
  SboxInst_n293 <= LPM_d0_ivl_6279(0);
  tmp_ivl_6282 <= y0(35);
  LPM_q_ivl_6284 <= new_AGEMA_signal_2599 & tmp_ivl_6282;
  new_AGEMA_signal_3075 <= LPM_d0_ivl_6286(1);
  SboxInst_n292 <= LPM_d0_ivl_6286(0);
  tmp_ivl_6289 <= y0(36);
  LPM_q_ivl_6291 <= new_AGEMA_signal_2597 & tmp_ivl_6289;
  new_AGEMA_signal_3076 <= LPM_d0_ivl_6293(1);
  SboxInst_n291 <= LPM_d0_ivl_6293(0);
  tmp_ivl_6296 <= y0(37);
  LPM_q_ivl_6298 <= new_AGEMA_signal_2595 & tmp_ivl_6296;
  new_AGEMA_signal_3077 <= LPM_d0_ivl_6300(1);
  SboxInst_n290 <= LPM_d0_ivl_6300(0);
  tmp_ivl_6303 <= y0(38);
  LPM_q_ivl_6305 <= new_AGEMA_signal_2593 & tmp_ivl_6303;
  new_AGEMA_signal_3078 <= LPM_d0_ivl_6307(1);
  SboxInst_n289 <= LPM_d0_ivl_6307(0);
  tmp_ivl_6310 <= y0(39);
  LPM_q_ivl_6312 <= new_AGEMA_signal_2591 & tmp_ivl_6310;
  new_AGEMA_signal_3079 <= LPM_d0_ivl_6314(1);
  SboxInst_n288 <= LPM_d0_ivl_6314(0);
  tmp_ivl_6317 <= y0(3);
  LPM_q_ivl_6319 <= new_AGEMA_signal_2589 & tmp_ivl_6317;
  new_AGEMA_signal_3080 <= LPM_d0_ivl_6321(1);
  SboxInst_n287 <= LPM_d0_ivl_6321(0);
  tmp_ivl_6324 <= y0(40);
  LPM_q_ivl_6326 <= new_AGEMA_signal_2587 & tmp_ivl_6324;
  new_AGEMA_signal_3081 <= LPM_d0_ivl_6328(1);
  SboxInst_n286 <= LPM_d0_ivl_6328(0);
  tmp_ivl_6331 <= y0(41);
  LPM_q_ivl_6333 <= new_AGEMA_signal_2585 & tmp_ivl_6331;
  new_AGEMA_signal_3082 <= LPM_d0_ivl_6335(1);
  SboxInst_n285 <= LPM_d0_ivl_6335(0);
  tmp_ivl_6338 <= y0(42);
  LPM_q_ivl_6340 <= new_AGEMA_signal_2583 & tmp_ivl_6338;
  new_AGEMA_signal_3083 <= LPM_d0_ivl_6342(1);
  SboxInst_n284 <= LPM_d0_ivl_6342(0);
  tmp_ivl_6345 <= y0(43);
  LPM_q_ivl_6347 <= new_AGEMA_signal_2581 & tmp_ivl_6345;
  new_AGEMA_signal_3084 <= LPM_d0_ivl_6349(1);
  SboxInst_n283 <= LPM_d0_ivl_6349(0);
  tmp_ivl_6352 <= y0(44);
  LPM_q_ivl_6354 <= new_AGEMA_signal_2579 & tmp_ivl_6352;
  new_AGEMA_signal_3085 <= LPM_d0_ivl_6356(1);
  SboxInst_n282 <= LPM_d0_ivl_6356(0);
  tmp_ivl_6359 <= y0(45);
  LPM_q_ivl_6361 <= new_AGEMA_signal_2577 & tmp_ivl_6359;
  new_AGEMA_signal_3086 <= LPM_d0_ivl_6363(1);
  SboxInst_n281 <= LPM_d0_ivl_6363(0);
  tmp_ivl_6366 <= y0(46);
  LPM_q_ivl_6368 <= new_AGEMA_signal_2575 & tmp_ivl_6366;
  new_AGEMA_signal_3087 <= LPM_d0_ivl_6370(1);
  SboxInst_n280 <= LPM_d0_ivl_6370(0);
  tmp_ivl_6373 <= y0(47);
  LPM_q_ivl_6375 <= new_AGEMA_signal_2573 & tmp_ivl_6373;
  new_AGEMA_signal_3088 <= LPM_d0_ivl_6377(1);
  SboxInst_n279 <= LPM_d0_ivl_6377(0);
  tmp_ivl_6380 <= y0(48);
  LPM_q_ivl_6382 <= new_AGEMA_signal_2571 & tmp_ivl_6380;
  new_AGEMA_signal_3089 <= LPM_d0_ivl_6384(1);
  SboxInst_n278 <= LPM_d0_ivl_6384(0);
  tmp_ivl_6387 <= y0(49);
  LPM_q_ivl_6389 <= new_AGEMA_signal_2569 & tmp_ivl_6387;
  new_AGEMA_signal_3090 <= LPM_d0_ivl_6391(1);
  SboxInst_n277 <= LPM_d0_ivl_6391(0);
  tmp_ivl_6394 <= y0(4);
  LPM_q_ivl_6396 <= new_AGEMA_signal_2567 & tmp_ivl_6394;
  new_AGEMA_signal_3091 <= LPM_d0_ivl_6398(1);
  SboxInst_n276 <= LPM_d0_ivl_6398(0);
  tmp_ivl_6401 <= y0(50);
  LPM_q_ivl_6403 <= new_AGEMA_signal_2565 & tmp_ivl_6401;
  new_AGEMA_signal_3092 <= LPM_d0_ivl_6405(1);
  SboxInst_n275 <= LPM_d0_ivl_6405(0);
  tmp_ivl_6408 <= y0(51);
  LPM_q_ivl_6410 <= new_AGEMA_signal_2563 & tmp_ivl_6408;
  new_AGEMA_signal_3093 <= LPM_d0_ivl_6412(1);
  SboxInst_n274 <= LPM_d0_ivl_6412(0);
  tmp_ivl_6415 <= y0(52);
  LPM_q_ivl_6417 <= new_AGEMA_signal_2561 & tmp_ivl_6415;
  new_AGEMA_signal_3094 <= LPM_d0_ivl_6419(1);
  SboxInst_n273 <= LPM_d0_ivl_6419(0);
  tmp_ivl_6422 <= y0(53);
  LPM_q_ivl_6424 <= new_AGEMA_signal_2559 & tmp_ivl_6422;
  new_AGEMA_signal_3095 <= LPM_d0_ivl_6426(1);
  SboxInst_n272 <= LPM_d0_ivl_6426(0);
  tmp_ivl_6429 <= y0(54);
  LPM_q_ivl_6431 <= new_AGEMA_signal_2557 & tmp_ivl_6429;
  new_AGEMA_signal_3096 <= LPM_d0_ivl_6433(1);
  SboxInst_n271 <= LPM_d0_ivl_6433(0);
  tmp_ivl_6436 <= y0(55);
  LPM_q_ivl_6438 <= new_AGEMA_signal_2555 & tmp_ivl_6436;
  new_AGEMA_signal_3097 <= LPM_d0_ivl_6440(1);
  SboxInst_n270 <= LPM_d0_ivl_6440(0);
  tmp_ivl_6443 <= y0(56);
  LPM_q_ivl_6445 <= new_AGEMA_signal_2553 & tmp_ivl_6443;
  new_AGEMA_signal_3098 <= LPM_d0_ivl_6447(1);
  SboxInst_n269 <= LPM_d0_ivl_6447(0);
  tmp_ivl_6450 <= y0(57);
  LPM_q_ivl_6452 <= new_AGEMA_signal_2551 & tmp_ivl_6450;
  new_AGEMA_signal_3099 <= LPM_d0_ivl_6454(1);
  SboxInst_n268 <= LPM_d0_ivl_6454(0);
  tmp_ivl_6457 <= y0(58);
  LPM_q_ivl_6459 <= new_AGEMA_signal_2549 & tmp_ivl_6457;
  new_AGEMA_signal_3100 <= LPM_d0_ivl_6461(1);
  SboxInst_n267 <= LPM_d0_ivl_6461(0);
  tmp_ivl_6464 <= y0(59);
  LPM_q_ivl_6466 <= new_AGEMA_signal_2547 & tmp_ivl_6464;
  new_AGEMA_signal_3101 <= LPM_d0_ivl_6468(1);
  SboxInst_n266 <= LPM_d0_ivl_6468(0);
  tmp_ivl_6471 <= y0(5);
  LPM_q_ivl_6473 <= new_AGEMA_signal_2545 & tmp_ivl_6471;
  new_AGEMA_signal_3102 <= LPM_d0_ivl_6475(1);
  SboxInst_n265 <= LPM_d0_ivl_6475(0);
  tmp_ivl_6478 <= y0(60);
  LPM_q_ivl_6480 <= new_AGEMA_signal_2543 & tmp_ivl_6478;
  new_AGEMA_signal_3103 <= LPM_d0_ivl_6482(1);
  SboxInst_n264 <= LPM_d0_ivl_6482(0);
  tmp_ivl_6485 <= y0(61);
  LPM_q_ivl_6487 <= new_AGEMA_signal_2541 & tmp_ivl_6485;
  new_AGEMA_signal_3104 <= LPM_d0_ivl_6489(1);
  SboxInst_n263 <= LPM_d0_ivl_6489(0);
  tmp_ivl_6492 <= y0(62);
  LPM_q_ivl_6494 <= new_AGEMA_signal_2539 & tmp_ivl_6492;
  new_AGEMA_signal_3105 <= LPM_d0_ivl_6496(1);
  SboxInst_n262 <= LPM_d0_ivl_6496(0);
  tmp_ivl_6499 <= y0(63);
  LPM_q_ivl_6501 <= new_AGEMA_signal_2537 & tmp_ivl_6499;
  new_AGEMA_signal_3106 <= LPM_d0_ivl_6503(1);
  SboxInst_n261 <= LPM_d0_ivl_6503(0);
  tmp_ivl_6506 <= y0(6);
  LPM_q_ivl_6508 <= new_AGEMA_signal_2535 & tmp_ivl_6506;
  new_AGEMA_signal_3107 <= LPM_d0_ivl_6510(1);
  SboxInst_n260 <= LPM_d0_ivl_6510(0);
  tmp_ivl_6513 <= y0(7);
  LPM_q_ivl_6515 <= new_AGEMA_signal_2533 & tmp_ivl_6513;
  new_AGEMA_signal_3108 <= LPM_d0_ivl_6517(1);
  SboxInst_n259 <= LPM_d0_ivl_6517(0);
  tmp_ivl_6520 <= y0(8);
  LPM_q_ivl_6522 <= new_AGEMA_signal_2531 & tmp_ivl_6520;
  new_AGEMA_signal_3109 <= LPM_d0_ivl_6524(1);
  SboxInst_n258 <= LPM_d0_ivl_6524(0);
  tmp_ivl_6527 <= y0(9);
  LPM_q_ivl_6529 <= new_AGEMA_signal_2529 & tmp_ivl_6527;
  new_AGEMA_signal_3110 <= LPM_d0_ivl_6531(1);
  SboxInst_n257 <= LPM_d0_ivl_6531(0);
  tmp_ivl_6534 <= state_in_s1(213);
  tmp_ivl_6536 <= state_in_s0(213);
  LPM_q_ivl_6538 <= tmp_ivl_6534 & tmp_ivl_6536;
  new_AGEMA_signal_2859 <= LPM_d0_ivl_6540(1);
  SboxInst_n345 <= LPM_d0_ivl_6540(0);
  tmp_ivl_6543 <= state_in_s1(223);
  tmp_ivl_6545 <= state_in_s0(223);
  LPM_q_ivl_6547 <= tmp_ivl_6543 & tmp_ivl_6545;
  new_AGEMA_signal_2860 <= LPM_d0_ivl_6549(1);
  SboxInst_n352 <= LPM_d0_ivl_6549(0);
  tmp_ivl_6552 <= state_in_s1(208);
  tmp_ivl_6554 <= state_in_s0(208);
  LPM_q_ivl_6556 <= tmp_ivl_6552 & tmp_ivl_6554;
  new_AGEMA_signal_2861 <= LPM_d0_ivl_6558(1);
  SboxInst_n350 <= LPM_d0_ivl_6558(0);
  tmp_ivl_6561 <= state_in_s1(212);
  tmp_ivl_6563 <= state_in_s0(212);
  LPM_q_ivl_6565 <= tmp_ivl_6561 & tmp_ivl_6563;
  new_AGEMA_signal_2862 <= LPM_d0_ivl_6567(1);
  SboxInst_n346 <= LPM_d0_ivl_6567(0);
  tmp_ivl_6570 <= state_in_s1(222);
  tmp_ivl_6572 <= state_in_s0(222);
  LPM_q_ivl_6574 <= tmp_ivl_6570 & tmp_ivl_6572;
  new_AGEMA_signal_2863 <= LPM_d0_ivl_6576(1);
  SboxInst_n353 <= LPM_d0_ivl_6576(0);
  tmp_ivl_6579 <= state_in_s1(211);
  tmp_ivl_6581 <= state_in_s0(211);
  LPM_q_ivl_6583 <= tmp_ivl_6579 & tmp_ivl_6581;
  new_AGEMA_signal_2864 <= LPM_d0_ivl_6585(1);
  SboxInst_n347 <= LPM_d0_ivl_6585(0);
  tmp_ivl_6588 <= state_in_s1(221);
  tmp_ivl_6590 <= state_in_s0(221);
  LPM_q_ivl_6592 <= tmp_ivl_6588 & tmp_ivl_6590;
  new_AGEMA_signal_2865 <= LPM_d0_ivl_6594(1);
  SboxInst_n354 <= LPM_d0_ivl_6594(0);
  tmp_ivl_6597 <= state_in_s1(210);
  tmp_ivl_6599 <= state_in_s0(210);
  LPM_q_ivl_6601 <= tmp_ivl_6597 & tmp_ivl_6599;
  new_AGEMA_signal_2866 <= LPM_d0_ivl_6603(1);
  SboxInst_n348 <= LPM_d0_ivl_6603(0);
  tmp_ivl_6606 <= state_in_s1(220);
  tmp_ivl_6608 <= state_in_s0(220);
  LPM_q_ivl_6610 <= tmp_ivl_6606 & tmp_ivl_6608;
  new_AGEMA_signal_2867 <= LPM_d0_ivl_6612(1);
  SboxInst_n355 <= LPM_d0_ivl_6612(0);
  tmp_ivl_6615 <= state_in_s1(209);
  tmp_ivl_6617 <= state_in_s0(209);
  LPM_q_ivl_6619 <= tmp_ivl_6615 & tmp_ivl_6617;
  new_AGEMA_signal_2868 <= LPM_d0_ivl_6621(1);
  SboxInst_n349 <= LPM_d0_ivl_6621(0);
  tmp_ivl_6624 <= state_in_s1(219);
  tmp_ivl_6626 <= state_in_s0(219);
  LPM_q_ivl_6628 <= tmp_ivl_6624 & tmp_ivl_6626;
  new_AGEMA_signal_2869 <= LPM_d0_ivl_6630(1);
  SboxInst_n356 <= LPM_d0_ivl_6630(0);
  tmp_ivl_6633 <= state_in_s1(218);
  tmp_ivl_6635 <= state_in_s0(218);
  LPM_q_ivl_6637 <= tmp_ivl_6633 & tmp_ivl_6635;
  new_AGEMA_signal_2870 <= LPM_d0_ivl_6639(1);
  SboxInst_n357 <= LPM_d0_ivl_6639(0);
  tmp_ivl_6642 <= state_in_s1(217);
  tmp_ivl_6644 <= state_in_s0(217);
  LPM_q_ivl_6646 <= tmp_ivl_6642 & tmp_ivl_6644;
  new_AGEMA_signal_2871 <= LPM_d0_ivl_6648(1);
  SboxInst_n358 <= LPM_d0_ivl_6648(0);
  tmp_ivl_6651 <= state_in_s1(216);
  tmp_ivl_6653 <= state_in_s0(216);
  LPM_q_ivl_6655 <= tmp_ivl_6651 & tmp_ivl_6653;
  new_AGEMA_signal_2872 <= LPM_d0_ivl_6657(1);
  SboxInst_n359 <= LPM_d0_ivl_6657(0);
  tmp_ivl_6660 <= state_in_s1(200);
  tmp_ivl_6662 <= state_in_s0(200);
  LPM_q_ivl_6664 <= tmp_ivl_6660 & tmp_ivl_6662;
  new_AGEMA_signal_2873 <= LPM_d0_ivl_6666(1);
  SboxInst_n342 <= LPM_d0_ivl_6666(0);
  tmp_ivl_6669 <= state_in_s1(205);
  tmp_ivl_6671 <= state_in_s0(205);
  LPM_q_ivl_6673 <= tmp_ivl_6669 & tmp_ivl_6671;
  new_AGEMA_signal_2874 <= LPM_d0_ivl_6675(1);
  SboxInst_n336 <= LPM_d0_ivl_6675(0);
  tmp_ivl_6678 <= state_in_s1(215);
  tmp_ivl_6680 <= state_in_s0(215);
  LPM_q_ivl_6682 <= tmp_ivl_6678 & tmp_ivl_6680;
  new_AGEMA_signal_2875 <= LPM_d0_ivl_6684(1);
  SboxInst_n343 <= LPM_d0_ivl_6684(0);
  tmp_ivl_6687 <= state_in_s1(204);
  tmp_ivl_6689 <= state_in_s0(204);
  LPM_q_ivl_6691 <= tmp_ivl_6687 & tmp_ivl_6689;
  new_AGEMA_signal_2876 <= LPM_d0_ivl_6693(1);
  SboxInst_n337 <= LPM_d0_ivl_6693(0);
  tmp_ivl_6696 <= state_in_s1(214);
  tmp_ivl_6698 <= state_in_s0(214);
  LPM_q_ivl_6700 <= tmp_ivl_6696 & tmp_ivl_6698;
  new_AGEMA_signal_2877 <= LPM_d0_ivl_6702(1);
  SboxInst_n344 <= LPM_d0_ivl_6702(0);
  tmp_ivl_6705 <= state_in_s1(203);
  tmp_ivl_6707 <= state_in_s0(203);
  LPM_q_ivl_6709 <= tmp_ivl_6705 & tmp_ivl_6707;
  new_AGEMA_signal_2878 <= LPM_d0_ivl_6711(1);
  SboxInst_n338 <= LPM_d0_ivl_6711(0);
  tmp_ivl_6714 <= state_in_s1(202);
  tmp_ivl_6716 <= state_in_s0(202);
  LPM_q_ivl_6718 <= tmp_ivl_6714 & tmp_ivl_6716;
  new_AGEMA_signal_2879 <= LPM_d0_ivl_6720(1);
  SboxInst_n339 <= LPM_d0_ivl_6720(0);
  tmp_ivl_6723 <= state_in_s1(201);
  tmp_ivl_6725 <= state_in_s0(201);
  LPM_q_ivl_6727 <= tmp_ivl_6723 & tmp_ivl_6725;
  new_AGEMA_signal_2880 <= LPM_d0_ivl_6729(1);
  SboxInst_n341 <= LPM_d0_ivl_6729(0);
  tmp_ivl_6732 <= state_in_s1(207);
  tmp_ivl_6734 <= state_in_s0(207);
  LPM_q_ivl_6736 <= tmp_ivl_6732 & tmp_ivl_6734;
  new_AGEMA_signal_2881 <= LPM_d0_ivl_6738(1);
  SboxInst_n334 <= LPM_d0_ivl_6738(0);
  tmp_ivl_6741 <= state_in_s1(197);
  tmp_ivl_6743 <= state_in_s0(197);
  LPM_q_ivl_6745 <= tmp_ivl_6741 & tmp_ivl_6743;
  new_AGEMA_signal_2882 <= LPM_d0_ivl_6747(1);
  SboxInst_n327 <= LPM_d0_ivl_6747(0);
  tmp_ivl_6750 <= state_in_s1(192);
  tmp_ivl_6752 <= state_in_s0(192);
  LPM_q_ivl_6754 <= tmp_ivl_6750 & tmp_ivl_6752;
  new_AGEMA_signal_2883 <= LPM_d0_ivl_6756(1);
  SboxInst_n333 <= LPM_d0_ivl_6756(0);
  tmp_ivl_6759 <= state_in_s1(206);
  tmp_ivl_6761 <= state_in_s0(206);
  LPM_q_ivl_6763 <= tmp_ivl_6759 & tmp_ivl_6761;
  new_AGEMA_signal_2884 <= LPM_d0_ivl_6765(1);
  SboxInst_n335 <= LPM_d0_ivl_6765(0);
  tmp_ivl_6768 <= state_in_s1(196);
  tmp_ivl_6770 <= state_in_s0(196);
  LPM_q_ivl_6772 <= tmp_ivl_6768 & tmp_ivl_6770;
  new_AGEMA_signal_2885 <= LPM_d0_ivl_6774(1);
  SboxInst_n328 <= LPM_d0_ivl_6774(0);
  tmp_ivl_6777 <= state_in_s1(195);
  tmp_ivl_6779 <= state_in_s0(195);
  LPM_q_ivl_6781 <= tmp_ivl_6777 & tmp_ivl_6779;
  new_AGEMA_signal_2886 <= LPM_d0_ivl_6783(1);
  SboxInst_n330 <= LPM_d0_ivl_6783(0);
  tmp_ivl_6786 <= state_in_s1(194);
  tmp_ivl_6788 <= state_in_s0(194);
  LPM_q_ivl_6790 <= tmp_ivl_6786 & tmp_ivl_6788;
  new_AGEMA_signal_2887 <= LPM_d0_ivl_6792(1);
  SboxInst_n331 <= LPM_d0_ivl_6792(0);
  tmp_ivl_6795 <= state_in_s1(193);
  tmp_ivl_6797 <= state_in_s0(193);
  LPM_q_ivl_6799 <= tmp_ivl_6795 & tmp_ivl_6797;
  new_AGEMA_signal_2888 <= LPM_d0_ivl_6801(1);
  SboxInst_n332 <= LPM_d0_ivl_6801(0);
  tmp_ivl_6804 <= state_in_s1(199);
  tmp_ivl_6806 <= state_in_s0(199);
  LPM_q_ivl_6808 <= tmp_ivl_6804 & tmp_ivl_6806;
  new_AGEMA_signal_2889 <= LPM_d0_ivl_6810(1);
  SboxInst_n325 <= LPM_d0_ivl_6810(0);
  tmp_ivl_6813 <= state_in_s1(248);
  tmp_ivl_6815 <= state_in_s0(248);
  LPM_q_ivl_6817 <= tmp_ivl_6813 & tmp_ivl_6815;
  new_AGEMA_signal_2890 <= LPM_d0_ivl_6819(1);
  SboxInst_n384 <= LPM_d0_ivl_6819(0);
  tmp_ivl_6822 <= state_in_s1(253);
  tmp_ivl_6824 <= state_in_s0(253);
  LPM_q_ivl_6826 <= tmp_ivl_6822 & tmp_ivl_6824;
  new_AGEMA_signal_2891 <= LPM_d0_ivl_6828(1);
  SboxInst_n329 <= LPM_d0_ivl_6828(0);
  tmp_ivl_6831 <= state_in_s1(252);
  tmp_ivl_6833 <= state_in_s0(252);
  LPM_q_ivl_6835 <= tmp_ivl_6831 & tmp_ivl_6833;
  new_AGEMA_signal_2892 <= LPM_d0_ivl_6837(1);
  SboxInst_n340 <= LPM_d0_ivl_6837(0);
  tmp_ivl_6840 <= state_in_s1(198);
  tmp_ivl_6842 <= state_in_s0(198);
  LPM_q_ivl_6844 <= tmp_ivl_6840 & tmp_ivl_6842;
  new_AGEMA_signal_2893 <= LPM_d0_ivl_6846(1);
  SboxInst_n326 <= LPM_d0_ivl_6846(0);
  tmp_ivl_6849 <= state_in_s1(251);
  tmp_ivl_6851 <= state_in_s0(251);
  LPM_q_ivl_6853 <= tmp_ivl_6849 & tmp_ivl_6851;
  new_AGEMA_signal_2894 <= LPM_d0_ivl_6855(1);
  SboxInst_n351 <= LPM_d0_ivl_6855(0);
  tmp_ivl_6858 <= state_in_s1(250);
  tmp_ivl_6860 <= state_in_s0(250);
  LPM_q_ivl_6862 <= tmp_ivl_6858 & tmp_ivl_6860;
  new_AGEMA_signal_2895 <= LPM_d0_ivl_6864(1);
  SboxInst_n362 <= LPM_d0_ivl_6864(0);
  tmp_ivl_6867 <= state_in_s1(249);
  tmp_ivl_6869 <= state_in_s0(249);
  LPM_q_ivl_6871 <= tmp_ivl_6867 & tmp_ivl_6869;
  new_AGEMA_signal_2896 <= LPM_d0_ivl_6873(1);
  SboxInst_n373 <= LPM_d0_ivl_6873(0);
  tmp_ivl_6876 <= state_in_s1(86);
  tmp_ivl_6878 <= state_in_s0(86);
  LPM_q_ivl_6880 <= tmp_ivl_6876 & tmp_ivl_6878;
  new_AGEMA_signal_2897 <= LPM_d0_ivl_6882(1);
  SboxInst_n216 <= LPM_d0_ivl_6882(0);
  tmp_ivl_6885 <= state_in_s1(127);
  tmp_ivl_6887 <= state_in_s0(127);
  LPM_q_ivl_6889 <= tmp_ivl_6885 & tmp_ivl_6887;
  new_AGEMA_signal_2899 <= LPM_d0_ivl_6891(1);
  SboxInst_n195 <= LPM_d0_ivl_6891(0);
  tmp_ivl_6894 <= state_in_s1(124);
  tmp_ivl_6896 <= state_in_s0(124);
  LPM_q_ivl_6898 <= tmp_ivl_6894 & tmp_ivl_6896;
  new_AGEMA_signal_2900 <= LPM_d0_ivl_6900(1);
  SboxInst_n212 <= LPM_d0_ivl_6900(0);
  tmp_ivl_6903 <= state_in_s1(126);
  tmp_ivl_6905 <= state_in_s0(126);
  LPM_q_ivl_6907 <= tmp_ivl_6903 & tmp_ivl_6905;
  new_AGEMA_signal_2901 <= LPM_d0_ivl_6909(1);
  SboxInst_n196 <= LPM_d0_ivl_6909(0);
  tmp_ivl_6912 <= state_in_s1(85);
  tmp_ivl_6914 <= state_in_s0(85);
  LPM_q_ivl_6916 <= tmp_ivl_6912 & tmp_ivl_6914;
  new_AGEMA_signal_2902 <= LPM_d0_ivl_6918(1);
  SboxInst_n217 <= LPM_d0_ivl_6918(0);
  tmp_ivl_6921 <= state_in_s1(123);
  tmp_ivl_6923 <= state_in_s0(123);
  LPM_q_ivl_6925 <= tmp_ivl_6921 & tmp_ivl_6923;
  new_AGEMA_signal_2904 <= LPM_d0_ivl_6927(1);
  SboxInst_n223 <= LPM_d0_ivl_6927(0);
  tmp_ivl_6930 <= state_in_s1(84);
  tmp_ivl_6932 <= state_in_s0(84);
  LPM_q_ivl_6934 <= tmp_ivl_6930 & tmp_ivl_6932;
  new_AGEMA_signal_2905 <= LPM_d0_ivl_6936(1);
  SboxInst_n218 <= LPM_d0_ivl_6936(0);
  tmp_ivl_6939 <= state_in_s1(122);
  tmp_ivl_6941 <= state_in_s0(122);
  LPM_q_ivl_6943 <= tmp_ivl_6939 & tmp_ivl_6941;
  new_AGEMA_signal_2906 <= LPM_d0_ivl_6945(1);
  SboxInst_n234 <= LPM_d0_ivl_6945(0);
  tmp_ivl_6948 <= state_in_s1(125);
  tmp_ivl_6950 <= state_in_s0(125);
  LPM_q_ivl_6952 <= tmp_ivl_6948 & tmp_ivl_6950;
  new_AGEMA_signal_2907 <= LPM_d0_ivl_6954(1);
  SboxInst_n201 <= LPM_d0_ivl_6954(0);
  tmp_ivl_6957 <= state_in_s1(83);
  tmp_ivl_6959 <= state_in_s0(83);
  LPM_q_ivl_6961 <= tmp_ivl_6957 & tmp_ivl_6959;
  new_AGEMA_signal_2908 <= LPM_d0_ivl_6963(1);
  SboxInst_n219 <= LPM_d0_ivl_6963(0);
  tmp_ivl_6966 <= state_in_s1(121);
  tmp_ivl_6968 <= state_in_s0(121);
  LPM_q_ivl_6970 <= tmp_ivl_6966 & tmp_ivl_6968;
  new_AGEMA_signal_2909 <= LPM_d0_ivl_6972(1);
  SboxInst_n245 <= LPM_d0_ivl_6972(0);
  tmp_ivl_6975 <= state_in_s1(82);
  tmp_ivl_6977 <= state_in_s0(82);
  LPM_q_ivl_6979 <= tmp_ivl_6975 & tmp_ivl_6977;
  new_AGEMA_signal_2910 <= LPM_d0_ivl_6981(1);
  SboxInst_n220 <= LPM_d0_ivl_6981(0);
  tmp_ivl_6984 <= state_in_s1(120);
  tmp_ivl_6986 <= state_in_s0(120);
  LPM_q_ivl_6988 <= tmp_ivl_6984 & tmp_ivl_6986;
  new_AGEMA_signal_2911 <= LPM_d0_ivl_6990(1);
  SboxInst_n256 <= LPM_d0_ivl_6990(0);
  tmp_ivl_6993 <= state_in_s1(71);
  tmp_ivl_6995 <= state_in_s0(71);
  LPM_q_ivl_6997 <= tmp_ivl_6993 & tmp_ivl_6995;
  new_AGEMA_signal_2912 <= LPM_d0_ivl_6999(1);
  SboxInst_n197 <= LPM_d0_ivl_6999(0);
  tmp_ivl_7002 <= state_in_s1(81);
  tmp_ivl_7004 <= state_in_s0(81);
  LPM_q_ivl_7006 <= tmp_ivl_7002 & tmp_ivl_7004;
  new_AGEMA_signal_2913 <= LPM_d0_ivl_7008(1);
  SboxInst_n221 <= LPM_d0_ivl_7008(0);
  tmp_ivl_7011 <= state_in_s1(80);
  tmp_ivl_7013 <= state_in_s0(80);
  LPM_q_ivl_7015 <= tmp_ivl_7011 & tmp_ivl_7013;
  new_AGEMA_signal_2914 <= LPM_d0_ivl_7017(1);
  SboxInst_n222 <= LPM_d0_ivl_7017(0);
  tmp_ivl_7020 <= state_in_s1(70);
  tmp_ivl_7022 <= state_in_s0(70);
  LPM_q_ivl_7024 <= tmp_ivl_7020 & tmp_ivl_7022;
  new_AGEMA_signal_2915 <= LPM_d0_ivl_7026(1);
  SboxInst_n198 <= LPM_d0_ivl_7026(0);
  tmp_ivl_7029 <= state_in_s1(95);
  tmp_ivl_7031 <= state_in_s0(95);
  LPM_q_ivl_7033 <= tmp_ivl_7029 & tmp_ivl_7031;
  new_AGEMA_signal_2916 <= LPM_d0_ivl_7035(1);
  SboxInst_n224 <= LPM_d0_ivl_7035(0);
  tmp_ivl_7038 <= state_in_s1(69);
  tmp_ivl_7040 <= state_in_s0(69);
  LPM_q_ivl_7042 <= tmp_ivl_7038 & tmp_ivl_7040;
  new_AGEMA_signal_2917 <= LPM_d0_ivl_7044(1);
  SboxInst_n199 <= LPM_d0_ivl_7044(0);
  tmp_ivl_7047 <= state_in_s1(119);
  tmp_ivl_7049 <= state_in_s0(119);
  LPM_q_ivl_7051 <= tmp_ivl_7047 & tmp_ivl_7049;
  new_AGEMA_signal_2918 <= LPM_d0_ivl_7053(1);
  SboxInst_n250 <= LPM_d0_ivl_7053(0);
  tmp_ivl_7056 <= state_in_s1(116);
  tmp_ivl_7058 <= state_in_s0(116);
  LPM_q_ivl_7060 <= tmp_ivl_7056 & tmp_ivl_7058;
  new_AGEMA_signal_2919 <= LPM_d0_ivl_7062(1);
  SboxInst_n253 <= LPM_d0_ivl_7062(0);
  tmp_ivl_7065 <= state_in_s1(78);
  tmp_ivl_7067 <= state_in_s0(78);
  LPM_q_ivl_7069 <= tmp_ivl_7065 & tmp_ivl_7067;
  new_AGEMA_signal_2920 <= LPM_d0_ivl_7071(1);
  SboxInst_n207 <= LPM_d0_ivl_7071(0);
  tmp_ivl_7074 <= state_in_s1(115);
  tmp_ivl_7076 <= state_in_s0(115);
  LPM_q_ivl_7078 <= tmp_ivl_7074 & tmp_ivl_7076;
  new_AGEMA_signal_2921 <= LPM_d0_ivl_7080(1);
  SboxInst_n254 <= LPM_d0_ivl_7080(0);
  tmp_ivl_7083 <= state_in_s1(118);
  tmp_ivl_7085 <= state_in_s0(118);
  LPM_q_ivl_7087 <= tmp_ivl_7083 & tmp_ivl_7085;
  new_AGEMA_signal_2922 <= LPM_d0_ivl_7089(1);
  SboxInst_n251 <= LPM_d0_ivl_7089(0);
  tmp_ivl_7092 <= state_in_s1(77);
  tmp_ivl_7094 <= state_in_s0(77);
  LPM_q_ivl_7096 <= tmp_ivl_7092 & tmp_ivl_7094;
  new_AGEMA_signal_2923 <= LPM_d0_ivl_7098(1);
  SboxInst_n208 <= LPM_d0_ivl_7098(0);
  tmp_ivl_7101 <= state_in_s1(114);
  tmp_ivl_7103 <= state_in_s0(114);
  LPM_q_ivl_7105 <= tmp_ivl_7101 & tmp_ivl_7103;
  new_AGEMA_signal_2924 <= LPM_d0_ivl_7107(1);
  SboxInst_n255 <= LPM_d0_ivl_7107(0);
  tmp_ivl_7110 <= state_in_s1(117);
  tmp_ivl_7112 <= state_in_s0(117);
  LPM_q_ivl_7114 <= tmp_ivl_7110 & tmp_ivl_7112;
  new_AGEMA_signal_2925 <= LPM_d0_ivl_7116(1);
  SboxInst_n252 <= LPM_d0_ivl_7116(0);
  tmp_ivl_7119 <= state_in_s1(76);
  tmp_ivl_7121 <= state_in_s0(76);
  LPM_q_ivl_7123 <= tmp_ivl_7119 & tmp_ivl_7121;
  new_AGEMA_signal_2926 <= LPM_d0_ivl_7125(1);
  SboxInst_n209 <= LPM_d0_ivl_7125(0);
  tmp_ivl_7128 <= state_in_s1(113);
  tmp_ivl_7130 <= state_in_s0(113);
  LPM_q_ivl_7132 <= tmp_ivl_7128 & tmp_ivl_7130;
  new_AGEMA_signal_2927 <= LPM_d0_ivl_7134(1);
  SboxInst_n193 <= LPM_d0_ivl_7134(0);
  tmp_ivl_7137 <= state_in_s1(75);
  tmp_ivl_7139 <= state_in_s0(75);
  LPM_q_ivl_7141 <= tmp_ivl_7137 & tmp_ivl_7139;
  new_AGEMA_signal_2928 <= LPM_d0_ivl_7143(1);
  SboxInst_n210 <= LPM_d0_ivl_7143(0);
  tmp_ivl_7146 <= state_in_s1(112);
  tmp_ivl_7148 <= state_in_s0(112);
  LPM_q_ivl_7150 <= tmp_ivl_7146 & tmp_ivl_7148;
  new_AGEMA_signal_2929 <= LPM_d0_ivl_7152(1);
  SboxInst_n194 <= LPM_d0_ivl_7152(0);
  tmp_ivl_7155 <= state_in_s1(74);
  tmp_ivl_7157 <= state_in_s0(74);
  LPM_q_ivl_7159 <= tmp_ivl_7155 & tmp_ivl_7157;
  new_AGEMA_signal_2930 <= LPM_d0_ivl_7161(1);
  SboxInst_n211 <= LPM_d0_ivl_7161(0);
  tmp_ivl_7164 <= state_in_s1(73);
  tmp_ivl_7166 <= state_in_s0(73);
  LPM_q_ivl_7168 <= tmp_ivl_7164 & tmp_ivl_7166;
  new_AGEMA_signal_2931 <= LPM_d0_ivl_7170(1);
  SboxInst_n213 <= LPM_d0_ivl_7170(0);
  tmp_ivl_7173 <= state_in_s1(72);
  tmp_ivl_7175 <= state_in_s0(72);
  LPM_q_ivl_7177 <= tmp_ivl_7173 & tmp_ivl_7175;
  new_AGEMA_signal_2932 <= LPM_d0_ivl_7179(1);
  SboxInst_n214 <= LPM_d0_ivl_7179(0);
  tmp_ivl_7182 <= state_in_s1(87);
  tmp_ivl_7184 <= state_in_s0(87);
  LPM_q_ivl_7186 <= tmp_ivl_7182 & tmp_ivl_7184;
  new_AGEMA_signal_2933 <= LPM_d0_ivl_7188(1);
  SboxInst_n215 <= LPM_d0_ivl_7188(0);
  tmp_ivl_7191 <= state_in_s1(108);
  tmp_ivl_7193 <= state_in_s0(108);
  LPM_q_ivl_7195 <= tmp_ivl_7191 & tmp_ivl_7193;
  new_AGEMA_signal_2934 <= LPM_d0_ivl_7197(1);
  SboxInst_n244 <= LPM_d0_ivl_7197(0);
  tmp_ivl_7200 <= state_in_s1(111);
  tmp_ivl_7202 <= state_in_s0(111);
  LPM_q_ivl_7204 <= tmp_ivl_7200 & tmp_ivl_7202;
  new_AGEMA_signal_2935 <= LPM_d0_ivl_7206(1);
  SboxInst_n241 <= LPM_d0_ivl_7206(0);
  tmp_ivl_7209 <= state_in_s1(107);
  tmp_ivl_7211 <= state_in_s0(107);
  LPM_q_ivl_7213 <= tmp_ivl_7209 & tmp_ivl_7211;
  new_AGEMA_signal_2936 <= LPM_d0_ivl_7215(1);
  SboxInst_n246 <= LPM_d0_ivl_7215(0);
  tmp_ivl_7218 <= state_in_s1(110);
  tmp_ivl_7220 <= state_in_s0(110);
  LPM_q_ivl_7222 <= tmp_ivl_7218 & tmp_ivl_7220;
  new_AGEMA_signal_2937 <= LPM_d0_ivl_7224(1);
  SboxInst_n242 <= LPM_d0_ivl_7224(0);
  tmp_ivl_7227 <= state_in_s1(68);
  tmp_ivl_7229 <= state_in_s0(68);
  LPM_q_ivl_7231 <= tmp_ivl_7227 & tmp_ivl_7229;
  new_AGEMA_signal_2938 <= LPM_d0_ivl_7233(1);
  SboxInst_n200 <= LPM_d0_ivl_7233(0);
  tmp_ivl_7236 <= state_in_s1(109);
  tmp_ivl_7238 <= state_in_s0(109);
  LPM_q_ivl_7240 <= tmp_ivl_7236 & tmp_ivl_7238;
  new_AGEMA_signal_2939 <= LPM_d0_ivl_7242(1);
  SboxInst_n243 <= LPM_d0_ivl_7242(0);
  tmp_ivl_7245 <= state_in_s1(106);
  tmp_ivl_7247 <= state_in_s0(106);
  LPM_q_ivl_7249 <= tmp_ivl_7245 & tmp_ivl_7247;
  new_AGEMA_signal_2940 <= LPM_d0_ivl_7251(1);
  SboxInst_n247 <= LPM_d0_ivl_7251(0);
  tmp_ivl_7254 <= state_in_s1(67);
  tmp_ivl_7256 <= state_in_s0(67);
  LPM_q_ivl_7258 <= tmp_ivl_7254 & tmp_ivl_7256;
  new_AGEMA_signal_2941 <= LPM_d0_ivl_7260(1);
  SboxInst_n202 <= LPM_d0_ivl_7260(0);
  tmp_ivl_7263 <= state_in_s1(105);
  tmp_ivl_7265 <= state_in_s0(105);
  LPM_q_ivl_7267 <= tmp_ivl_7263 & tmp_ivl_7265;
  new_AGEMA_signal_2942 <= LPM_d0_ivl_7269(1);
  SboxInst_n248 <= LPM_d0_ivl_7269(0);
  tmp_ivl_7272 <= state_in_s1(66);
  tmp_ivl_7274 <= state_in_s0(66);
  LPM_q_ivl_7276 <= tmp_ivl_7272 & tmp_ivl_7274;
  new_AGEMA_signal_2943 <= LPM_d0_ivl_7278(1);
  SboxInst_n203 <= LPM_d0_ivl_7278(0);
  tmp_ivl_7281 <= state_in_s1(104);
  tmp_ivl_7283 <= state_in_s0(104);
  LPM_q_ivl_7285 <= tmp_ivl_7281 & tmp_ivl_7283;
  new_AGEMA_signal_2944 <= LPM_d0_ivl_7287(1);
  SboxInst_n249 <= LPM_d0_ivl_7287(0);
  tmp_ivl_7290 <= state_in_s1(65);
  tmp_ivl_7292 <= state_in_s0(65);
  LPM_q_ivl_7294 <= tmp_ivl_7290 & tmp_ivl_7292;
  new_AGEMA_signal_2945 <= LPM_d0_ivl_7296(1);
  SboxInst_n204 <= LPM_d0_ivl_7296(0);
  tmp_ivl_7299 <= state_in_s1(64);
  tmp_ivl_7301 <= state_in_s0(64);
  LPM_q_ivl_7303 <= tmp_ivl_7299 & tmp_ivl_7301;
  new_AGEMA_signal_2946 <= LPM_d0_ivl_7305(1);
  SboxInst_n205 <= LPM_d0_ivl_7305(0);
  tmp_ivl_7308 <= state_in_s1(79);
  tmp_ivl_7310 <= state_in_s0(79);
  LPM_q_ivl_7312 <= tmp_ivl_7308 & tmp_ivl_7310;
  new_AGEMA_signal_2947 <= LPM_d0_ivl_7314(1);
  SboxInst_n206 <= LPM_d0_ivl_7314(0);
  tmp_ivl_7317 <= state_in_s1(103);
  tmp_ivl_7319 <= state_in_s0(103);
  LPM_q_ivl_7321 <= tmp_ivl_7317 & tmp_ivl_7319;
  new_AGEMA_signal_2948 <= LPM_d0_ivl_7323(1);
  SboxInst_n232 <= LPM_d0_ivl_7323(0);
  tmp_ivl_7326 <= state_in_s1(100);
  tmp_ivl_7328 <= state_in_s0(100);
  LPM_q_ivl_7330 <= tmp_ivl_7326 & tmp_ivl_7328;
  new_AGEMA_signal_2949 <= LPM_d0_ivl_7332(1);
  SboxInst_n236 <= LPM_d0_ivl_7332(0);
  tmp_ivl_7335 <= state_in_s1(102);
  tmp_ivl_7337 <= state_in_s0(102);
  LPM_q_ivl_7339 <= tmp_ivl_7335 & tmp_ivl_7337;
  new_AGEMA_signal_2950 <= LPM_d0_ivl_7341(1);
  SboxInst_n233 <= LPM_d0_ivl_7341(0);
  tmp_ivl_7344 <= state_in_s1(99);
  tmp_ivl_7346 <= state_in_s0(99);
  LPM_q_ivl_7348 <= tmp_ivl_7344 & tmp_ivl_7346;
  new_AGEMA_signal_2951 <= LPM_d0_ivl_7350(1);
  SboxInst_n237 <= LPM_d0_ivl_7350(0);
  tmp_ivl_7353 <= state_in_s1(98);
  tmp_ivl_7355 <= state_in_s0(98);
  LPM_q_ivl_7357 <= tmp_ivl_7353 & tmp_ivl_7355;
  new_AGEMA_signal_2952 <= LPM_d0_ivl_7359(1);
  SboxInst_n238 <= LPM_d0_ivl_7359(0);
  tmp_ivl_7362 <= state_in_s1(101);
  tmp_ivl_7364 <= state_in_s0(101);
  LPM_q_ivl_7366 <= tmp_ivl_7362 & tmp_ivl_7364;
  new_AGEMA_signal_2953 <= LPM_d0_ivl_7368(1);
  SboxInst_n235 <= LPM_d0_ivl_7368(0);
  tmp_ivl_7371 <= state_in_s1(97);
  tmp_ivl_7373 <= state_in_s0(97);
  LPM_q_ivl_7375 <= tmp_ivl_7371 & tmp_ivl_7373;
  new_AGEMA_signal_2954 <= LPM_d0_ivl_7377(1);
  SboxInst_n239 <= LPM_d0_ivl_7377(0);
  tmp_ivl_7380 <= state_in_s1(96);
  tmp_ivl_7382 <= state_in_s0(96);
  LPM_q_ivl_7384 <= tmp_ivl_7380 & tmp_ivl_7382;
  new_AGEMA_signal_2955 <= LPM_d0_ivl_7386(1);
  SboxInst_n240 <= LPM_d0_ivl_7386(0);
  tmp_ivl_7389 <= state_in_s1(92);
  tmp_ivl_7391 <= state_in_s0(92);
  LPM_q_ivl_7393 <= tmp_ivl_7389 & tmp_ivl_7391;
  new_AGEMA_signal_2956 <= LPM_d0_ivl_7395(1);
  SboxInst_n227 <= LPM_d0_ivl_7395(0);
  tmp_ivl_7398 <= state_in_s1(91);
  tmp_ivl_7400 <= state_in_s0(91);
  LPM_q_ivl_7402 <= tmp_ivl_7398 & tmp_ivl_7400;
  new_AGEMA_signal_2957 <= LPM_d0_ivl_7404(1);
  SboxInst_n228 <= LPM_d0_ivl_7404(0);
  tmp_ivl_7407 <= state_in_s1(94);
  tmp_ivl_7409 <= state_in_s0(94);
  LPM_q_ivl_7411 <= tmp_ivl_7407 & tmp_ivl_7409;
  new_AGEMA_signal_2958 <= LPM_d0_ivl_7413(1);
  SboxInst_n225 <= LPM_d0_ivl_7413(0);
  tmp_ivl_7416 <= state_in_s1(90);
  tmp_ivl_7418 <= state_in_s0(90);
  LPM_q_ivl_7420 <= tmp_ivl_7416 & tmp_ivl_7418;
  new_AGEMA_signal_2959 <= LPM_d0_ivl_7422(1);
  SboxInst_n229 <= LPM_d0_ivl_7422(0);
  tmp_ivl_7425 <= state_in_s1(93);
  tmp_ivl_7427 <= state_in_s0(93);
  LPM_q_ivl_7429 <= tmp_ivl_7425 & tmp_ivl_7427;
  new_AGEMA_signal_2960 <= LPM_d0_ivl_7431(1);
  SboxInst_n226 <= LPM_d0_ivl_7431(0);
  tmp_ivl_7434 <= state_in_s1(89);
  tmp_ivl_7436 <= state_in_s0(89);
  LPM_q_ivl_7438 <= tmp_ivl_7434 & tmp_ivl_7436;
  new_AGEMA_signal_2961 <= LPM_d0_ivl_7440(1);
  SboxInst_n230 <= LPM_d0_ivl_7440(0);
  tmp_ivl_7443 <= state_in_s1(88);
  tmp_ivl_7445 <= state_in_s0(88);
  LPM_q_ivl_7447 <= tmp_ivl_7443 & tmp_ivl_7445;
  new_AGEMA_signal_2962 <= LPM_d0_ivl_7449(1);
  SboxInst_n231 <= LPM_d0_ivl_7449(0);
  tmp_ivl_7452 <= state_in_s1(255);
  tmp_ivl_7454 <= state_in_s0(255);
  LPM_q_ivl_7456 <= tmp_ivl_7452 & tmp_ivl_7454;
  new_AGEMA_signal_2963 <= LPM_d0_ivl_7458(1);
  SboxInst_n323 <= LPM_d0_ivl_7458(0);
  tmp_ivl_7461 <= state_in_s1(233);
  tmp_ivl_7463 <= state_in_s0(233);
  LPM_q_ivl_7465 <= tmp_ivl_7461 & tmp_ivl_7463;
  new_AGEMA_signal_2964 <= LPM_d0_ivl_7467(1);
  SboxInst_n376 <= LPM_d0_ivl_7467(0);
  tmp_ivl_7470 <= state_in_s1(224);
  tmp_ivl_7472 <= state_in_s0(224);
  LPM_q_ivl_7474 <= tmp_ivl_7470 & tmp_ivl_7472;
  new_AGEMA_signal_2965 <= LPM_d0_ivl_7476(1);
  SboxInst_n368 <= LPM_d0_ivl_7476(0);
  tmp_ivl_7479 <= state_in_s1(254);
  tmp_ivl_7481 <= state_in_s0(254);
  LPM_q_ivl_7483 <= tmp_ivl_7479 & tmp_ivl_7481;
  new_AGEMA_signal_2966 <= LPM_d0_ivl_7485(1);
  SboxInst_n324 <= LPM_d0_ivl_7485(0);
  tmp_ivl_7488 <= state_in_s1(239);
  tmp_ivl_7490 <= state_in_s0(239);
  LPM_q_ivl_7492 <= tmp_ivl_7488 & tmp_ivl_7490;
  new_AGEMA_signal_2967 <= LPM_d0_ivl_7494(1);
  SboxInst_n369 <= LPM_d0_ivl_7494(0);
  tmp_ivl_7497 <= state_in_s1(232);
  tmp_ivl_7499 <= state_in_s0(232);
  LPM_q_ivl_7501 <= tmp_ivl_7497 & tmp_ivl_7499;
  new_AGEMA_signal_2968 <= LPM_d0_ivl_7503(1);
  SboxInst_n377 <= LPM_d0_ivl_7503(0);
  tmp_ivl_7506 <= state_in_s1(238);
  tmp_ivl_7508 <= state_in_s0(238);
  LPM_q_ivl_7510 <= tmp_ivl_7506 & tmp_ivl_7508;
  new_AGEMA_signal_2969 <= LPM_d0_ivl_7512(1);
  SboxInst_n370 <= LPM_d0_ivl_7512(0);
  tmp_ivl_7515 <= state_in_s1(247);
  tmp_ivl_7517 <= state_in_s0(247);
  LPM_q_ivl_7519 <= tmp_ivl_7515 & tmp_ivl_7517;
  new_AGEMA_signal_2970 <= LPM_d0_ivl_7521(1);
  SboxInst_n378 <= LPM_d0_ivl_7521(0);
  tmp_ivl_7524 <= state_in_s1(246);
  tmp_ivl_7526 <= state_in_s0(246);
  LPM_q_ivl_7528 <= tmp_ivl_7524 & tmp_ivl_7526;
  new_AGEMA_signal_2971 <= LPM_d0_ivl_7530(1);
  SboxInst_n379 <= LPM_d0_ivl_7530(0);
  tmp_ivl_7533 <= state_in_s1(237);
  tmp_ivl_7535 <= state_in_s0(237);
  LPM_q_ivl_7537 <= tmp_ivl_7533 & tmp_ivl_7535;
  new_AGEMA_signal_2972 <= LPM_d0_ivl_7539(1);
  SboxInst_n371 <= LPM_d0_ivl_7539(0);
  tmp_ivl_7542 <= state_in_s1(236);
  tmp_ivl_7544 <= state_in_s0(236);
  LPM_q_ivl_7546 <= tmp_ivl_7542 & tmp_ivl_7544;
  new_AGEMA_signal_2973 <= LPM_d0_ivl_7548(1);
  SboxInst_n372 <= LPM_d0_ivl_7548(0);
  tmp_ivl_7551 <= state_in_s1(245);
  tmp_ivl_7553 <= state_in_s0(245);
  LPM_q_ivl_7555 <= tmp_ivl_7551 & tmp_ivl_7553;
  new_AGEMA_signal_2974 <= LPM_d0_ivl_7557(1);
  SboxInst_n380 <= LPM_d0_ivl_7557(0);
  tmp_ivl_7560 <= state_in_s1(244);
  tmp_ivl_7562 <= state_in_s0(244);
  LPM_q_ivl_7564 <= tmp_ivl_7560 & tmp_ivl_7562;
  new_AGEMA_signal_2975 <= LPM_d0_ivl_7566(1);
  SboxInst_n381 <= LPM_d0_ivl_7566(0);
  tmp_ivl_7569 <= state_in_s1(235);
  tmp_ivl_7571 <= state_in_s0(235);
  LPM_q_ivl_7573 <= tmp_ivl_7569 & tmp_ivl_7571;
  new_AGEMA_signal_2976 <= LPM_d0_ivl_7575(1);
  SboxInst_n374 <= LPM_d0_ivl_7575(0);
  tmp_ivl_7578 <= state_in_s1(243);
  tmp_ivl_7580 <= state_in_s0(243);
  LPM_q_ivl_7582 <= tmp_ivl_7578 & tmp_ivl_7580;
  new_AGEMA_signal_2977 <= LPM_d0_ivl_7584(1);
  SboxInst_n382 <= LPM_d0_ivl_7584(0);
  tmp_ivl_7587 <= state_in_s1(234);
  tmp_ivl_7589 <= state_in_s0(234);
  LPM_q_ivl_7591 <= tmp_ivl_7587 & tmp_ivl_7589;
  new_AGEMA_signal_2978 <= LPM_d0_ivl_7593(1);
  SboxInst_n375 <= LPM_d0_ivl_7593(0);
  tmp_ivl_7596 <= state_in_s1(242);
  tmp_ivl_7598 <= state_in_s0(242);
  LPM_q_ivl_7600 <= tmp_ivl_7596 & tmp_ivl_7598;
  new_AGEMA_signal_2979 <= LPM_d0_ivl_7602(1);
  SboxInst_n383 <= LPM_d0_ivl_7602(0);
  tmp_ivl_7605 <= state_in_s1(225);
  tmp_ivl_7607 <= state_in_s0(225);
  LPM_q_ivl_7609 <= tmp_ivl_7605 & tmp_ivl_7607;
  new_AGEMA_signal_2980 <= LPM_d0_ivl_7611(1);
  SboxInst_n367 <= LPM_d0_ivl_7611(0);
  tmp_ivl_7614 <= state_in_s1(231);
  tmp_ivl_7616 <= state_in_s0(231);
  LPM_q_ivl_7618 <= tmp_ivl_7614 & tmp_ivl_7616;
  new_AGEMA_signal_2981 <= LPM_d0_ivl_7620(1);
  SboxInst_n360 <= LPM_d0_ivl_7620(0);
  tmp_ivl_7623 <= state_in_s1(230);
  tmp_ivl_7625 <= state_in_s0(230);
  LPM_q_ivl_7627 <= tmp_ivl_7623 & tmp_ivl_7625;
  new_AGEMA_signal_2982 <= LPM_d0_ivl_7629(1);
  SboxInst_n361 <= LPM_d0_ivl_7629(0);
  tmp_ivl_7632 <= state_in_s1(229);
  tmp_ivl_7634 <= state_in_s0(229);
  LPM_q_ivl_7636 <= tmp_ivl_7632 & tmp_ivl_7634;
  new_AGEMA_signal_2983 <= LPM_d0_ivl_7638(1);
  SboxInst_n363 <= LPM_d0_ivl_7638(0);
  tmp_ivl_7641 <= state_in_s1(228);
  tmp_ivl_7643 <= state_in_s0(228);
  LPM_q_ivl_7645 <= tmp_ivl_7641 & tmp_ivl_7643;
  new_AGEMA_signal_2984 <= LPM_d0_ivl_7647(1);
  SboxInst_n364 <= LPM_d0_ivl_7647(0);
  tmp_ivl_7650 <= state_in_s1(227);
  tmp_ivl_7652 <= state_in_s0(227);
  LPM_q_ivl_7654 <= tmp_ivl_7650 & tmp_ivl_7652;
  new_AGEMA_signal_2985 <= LPM_d0_ivl_7656(1);
  SboxInst_n365 <= LPM_d0_ivl_7656(0);
  tmp_ivl_7659 <= state_in_s1(241);
  tmp_ivl_7661 <= state_in_s0(241);
  LPM_q_ivl_7663 <= tmp_ivl_7659 & tmp_ivl_7661;
  new_AGEMA_signal_2986 <= LPM_d0_ivl_7665(1);
  SboxInst_n321 <= LPM_d0_ivl_7665(0);
  tmp_ivl_7668 <= state_in_s1(226);
  tmp_ivl_7670 <= state_in_s0(226);
  LPM_q_ivl_7672 <= tmp_ivl_7668 & tmp_ivl_7670;
  new_AGEMA_signal_2987 <= LPM_d0_ivl_7674(1);
  SboxInst_n366 <= LPM_d0_ivl_7674(0);
  tmp_ivl_7677 <= state_in_s1(240);
  tmp_ivl_7679 <= state_in_s0(240);
  LPM_q_ivl_7681 <= tmp_ivl_7677 & tmp_ivl_7679;
  new_AGEMA_signal_2988 <= LPM_d0_ivl_7683(1);
  SboxInst_n322 <= LPM_d0_ivl_7683(0);
  tmp_ivl_7686 <= state_in_s1(238);
  tmp_ivl_7688 <= state_in_s0(238);
  tmp_ivl_7689 <= tmp_ivl_7686 & tmp_ivl_7688;
  LPM_q_ivl_7692 <= tmp_ivl_7694 & tmp_ivl_7689;
  tmp_ivl_7697 <= z4(22);
  tmp_ivl_7698 <= new_AGEMA_signal_3125 & tmp_ivl_7697;
  LPM_q_ivl_7701 <= tmp_ivl_7703 & tmp_ivl_7698;
  new_AGEMA_signal_3295 <= tmp_ivl_7705(1);
  n3405 <= tmp_ivl_7705(0);
  tmp_ivl_7705 <= LPM_d0_ivl_7709(0 + 1 downto 0);
  tmp_ivl_7711 <= state_in_s1(302);
  tmp_ivl_7713 <= state_in_s0(302);
  tmp_ivl_7714 <= tmp_ivl_7711 & tmp_ivl_7713;
  LPM_q_ivl_7717 <= tmp_ivl_7719 & tmp_ivl_7714;
  tmp_ivl_7721 <= new_AGEMA_signal_3295 & n3405;
  LPM_q_ivl_7724 <= tmp_ivl_7726 & tmp_ivl_7721;
  new_AGEMA_signal_3585 <= tmp_ivl_7728(1);
  n3926 <= tmp_ivl_7728(0);
  tmp_ivl_7728 <= LPM_d0_ivl_7732(0 + 1 downto 0);
  tmp_ivl_7734 <= state_in_s1(247);
  tmp_ivl_7736 <= state_in_s0(247);
  tmp_ivl_7737 <= tmp_ivl_7734 & tmp_ivl_7736;
  LPM_q_ivl_7740 <= tmp_ivl_7742 & tmp_ivl_7737;
  tmp_ivl_7745 <= z4(15);
  tmp_ivl_7746 <= new_AGEMA_signal_3117 & tmp_ivl_7745;
  LPM_q_ivl_7749 <= tmp_ivl_7751 & tmp_ivl_7746;
  new_AGEMA_signal_3296 <= tmp_ivl_7753(1);
  n3487 <= tmp_ivl_7753(0);
  tmp_ivl_7753 <= LPM_d0_ivl_7757(0 + 1 downto 0);
  tmp_ivl_7759 <= state_in_s1(311);
  tmp_ivl_7761 <= state_in_s0(311);
  tmp_ivl_7762 <= tmp_ivl_7759 & tmp_ivl_7761;
  LPM_q_ivl_7765 <= tmp_ivl_7767 & tmp_ivl_7762;
  tmp_ivl_7769 <= new_AGEMA_signal_3296 & n3487;
  LPM_q_ivl_7772 <= tmp_ivl_7774 & tmp_ivl_7769;
  new_AGEMA_signal_3586 <= tmp_ivl_7776(1);
  n3664 <= tmp_ivl_7776(0);
  tmp_ivl_7776 <= LPM_d0_ivl_7780(0 + 1 downto 0);
  tmp_ivl_7781 <= new_AGEMA_signal_3585 & n3926;
  LPM_q_ivl_7784 <= tmp_ivl_7786 & tmp_ivl_7781;
  tmp_ivl_7788 <= new_AGEMA_signal_3586 & n3664;
  LPM_q_ivl_7791 <= tmp_ivl_7793 & tmp_ivl_7788;
  new_AGEMA_signal_3891 <= tmp_ivl_7795(1);
  n3292 <= tmp_ivl_7795(0);
  tmp_ivl_7795 <= LPM_d0_ivl_7799(0 + 1 downto 0);
  tmp_ivl_7801 <= state_in_s1(192);
  tmp_ivl_7803 <= state_in_s0(192);
  tmp_ivl_7804 <= tmp_ivl_7801 & tmp_ivl_7803;
  LPM_q_ivl_7807 <= tmp_ivl_7809 & tmp_ivl_7804;
  tmp_ivl_7812 <= z4(56);
  tmp_ivl_7813 <= new_AGEMA_signal_3162 & tmp_ivl_7812;
  LPM_q_ivl_7816 <= tmp_ivl_7818 & tmp_ivl_7813;
  new_AGEMA_signal_3297 <= tmp_ivl_7820(1);
  n3441 <= tmp_ivl_7820(0);
  tmp_ivl_7820 <= LPM_d0_ivl_7824(0 + 1 downto 0);
  tmp_ivl_7826 <= state_in_s1(256);
  tmp_ivl_7828 <= state_in_s0(256);
  tmp_ivl_7829 <= tmp_ivl_7826 & tmp_ivl_7828;
  LPM_q_ivl_7832 <= tmp_ivl_7834 & tmp_ivl_7829;
  tmp_ivl_7836 <= new_AGEMA_signal_3297 & n3441;
  LPM_q_ivl_7839 <= tmp_ivl_7841 & tmp_ivl_7836;
  new_AGEMA_signal_3587 <= tmp_ivl_7843(1);
  n3657 <= tmp_ivl_7843(0);
  tmp_ivl_7843 <= LPM_d0_ivl_7847(0 + 1 downto 0);
  tmp_ivl_7848 <= new_AGEMA_signal_3891 & n3292;
  LPM_q_ivl_7851 <= tmp_ivl_7853 & tmp_ivl_7848;
  tmp_ivl_7855 <= new_AGEMA_signal_3587 & n3657;
  LPM_q_ivl_7858 <= tmp_ivl_7860 & tmp_ivl_7855;
  tmp_ivl_7862 <= tmp_ivl_7866(1);
  tmp_ivl_7864 <= tmp_ivl_7866(0);
  tmp_ivl_7866 <= LPM_d0_ivl_7870(0 + 1 downto 0);
  tmp_ivl_7872 <= state_in_s1(240);
  tmp_ivl_7874 <= state_in_s0(240);
  tmp_ivl_7875 <= tmp_ivl_7872 & tmp_ivl_7874;
  LPM_q_ivl_7878 <= tmp_ivl_7880 & tmp_ivl_7875;
  tmp_ivl_7883 <= z4(8);
  tmp_ivl_7884 <= new_AGEMA_signal_3173 & tmp_ivl_7883;
  LPM_q_ivl_7887 <= tmp_ivl_7889 & tmp_ivl_7884;
  new_AGEMA_signal_3298 <= tmp_ivl_7891(1);
  n3419 <= tmp_ivl_7891(0);
  tmp_ivl_7891 <= LPM_d0_ivl_7895(0 + 1 downto 0);
  tmp_ivl_7897 <= state_in_s1(304);
  tmp_ivl_7899 <= state_in_s0(304);
  tmp_ivl_7900 <= tmp_ivl_7897 & tmp_ivl_7899;
  LPM_q_ivl_7903 <= tmp_ivl_7905 & tmp_ivl_7900;
  tmp_ivl_7907 <= new_AGEMA_signal_3298 & n3419;
  LPM_q_ivl_7910 <= tmp_ivl_7912 & tmp_ivl_7907;
  new_AGEMA_signal_3588 <= tmp_ivl_7914(1);
  n3663 <= tmp_ivl_7914(0);
  tmp_ivl_7914 <= LPM_d0_ivl_7918(0 + 1 downto 0);
  tmp_ivl_7920 <= state_in_s1(210);
  tmp_ivl_7922 <= state_in_s0(210);
  tmp_ivl_7923 <= tmp_ivl_7920 & tmp_ivl_7922;
  LPM_q_ivl_7926 <= tmp_ivl_7928 & tmp_ivl_7923;
  tmp_ivl_7931 <= z4(42);
  tmp_ivl_7932 <= new_AGEMA_signal_3147 & tmp_ivl_7931;
  LPM_q_ivl_7935 <= tmp_ivl_7937 & tmp_ivl_7932;
  new_AGEMA_signal_3299 <= tmp_ivl_7939(1);
  n3615 <= tmp_ivl_7939(0);
  tmp_ivl_7939 <= LPM_d0_ivl_7943(0 + 1 downto 0);
  tmp_ivl_7945 <= state_in_s1(274);
  tmp_ivl_7947 <= state_in_s0(274);
  tmp_ivl_7948 <= tmp_ivl_7945 & tmp_ivl_7947;
  LPM_q_ivl_7951 <= tmp_ivl_7953 & tmp_ivl_7948;
  tmp_ivl_7955 <= new_AGEMA_signal_3299 & n3615;
  LPM_q_ivl_7958 <= tmp_ivl_7960 & tmp_ivl_7955;
  new_AGEMA_signal_3589 <= tmp_ivl_7962(1);
  n3661 <= tmp_ivl_7962(0);
  tmp_ivl_7962 <= LPM_d0_ivl_7966(0 + 1 downto 0);
  tmp_ivl_7967 <= new_AGEMA_signal_3588 & n3663;
  LPM_q_ivl_7970 <= tmp_ivl_7972 & tmp_ivl_7967;
  tmp_ivl_7974 <= new_AGEMA_signal_3589 & n3661;
  LPM_q_ivl_7977 <= tmp_ivl_7979 & tmp_ivl_7974;
  new_AGEMA_signal_3892 <= tmp_ivl_7981(1);
  n3293 <= tmp_ivl_7981(0);
  tmp_ivl_7981 <= LPM_d0_ivl_7985(0 + 1 downto 0);
  tmp_ivl_7987 <= state_in_s1(249);
  tmp_ivl_7989 <= state_in_s0(249);
  tmp_ivl_7990 <= tmp_ivl_7987 & tmp_ivl_7989;
  LPM_q_ivl_7993 <= tmp_ivl_7995 & tmp_ivl_7990;
  tmp_ivl_7998 <= z4(1);
  tmp_ivl_7999 <= new_AGEMA_signal_3122 & tmp_ivl_7998;
  LPM_q_ivl_8002 <= tmp_ivl_8004 & tmp_ivl_7999;
  new_AGEMA_signal_3300 <= tmp_ivl_8006(1);
  n3668 <= tmp_ivl_8006(0);
  tmp_ivl_8006 <= LPM_d0_ivl_8010(0 + 1 downto 0);
  tmp_ivl_8012 <= state_in_s1(313);
  tmp_ivl_8014 <= state_in_s0(313);
  tmp_ivl_8015 <= tmp_ivl_8012 & tmp_ivl_8014;
  LPM_q_ivl_8018 <= tmp_ivl_8020 & tmp_ivl_8015;
  tmp_ivl_8022 <= new_AGEMA_signal_3300 & n3668;
  LPM_q_ivl_8025 <= tmp_ivl_8027 & tmp_ivl_8022;
  new_AGEMA_signal_3590 <= tmp_ivl_8029(1);
  n3351 <= tmp_ivl_8029(0);
  tmp_ivl_8029 <= LPM_d0_ivl_8033(0 + 1 downto 0);
  tmp_ivl_8034 <= new_AGEMA_signal_3892 & n3293;
  LPM_q_ivl_8037 <= tmp_ivl_8039 & tmp_ivl_8034;
  tmp_ivl_8041 <= new_AGEMA_signal_3590 & n3351;
  LPM_q_ivl_8044 <= tmp_ivl_8046 & tmp_ivl_8041;
  tmp_ivl_8048 <= tmp_ivl_8052(1);
  tmp_ivl_8050 <= tmp_ivl_8052(0);
  tmp_ivl_8052 <= LPM_d0_ivl_8056(0 + 1 downto 0);
  tmp_ivl_8058 <= state_in_s1(241);
  tmp_ivl_8060 <= state_in_s0(241);
  tmp_ivl_8061 <= tmp_ivl_8058 & tmp_ivl_8060;
  LPM_q_ivl_8064 <= tmp_ivl_8066 & tmp_ivl_8061;
  tmp_ivl_8069 <= z4(9);
  tmp_ivl_8070 <= new_AGEMA_signal_3174 & tmp_ivl_8069;
  LPM_q_ivl_8073 <= tmp_ivl_8075 & tmp_ivl_8070;
  new_AGEMA_signal_3301 <= tmp_ivl_8077(1);
  n3478 <= tmp_ivl_8077(0);
  tmp_ivl_8077 <= LPM_d0_ivl_8081(0 + 1 downto 0);
  tmp_ivl_8083 <= state_in_s1(305);
  tmp_ivl_8085 <= state_in_s0(305);
  tmp_ivl_8086 <= tmp_ivl_8083 & tmp_ivl_8085;
  LPM_q_ivl_8089 <= tmp_ivl_8091 & tmp_ivl_8086;
  tmp_ivl_8093 <= new_AGEMA_signal_3301 & n3478;
  LPM_q_ivl_8096 <= tmp_ivl_8098 & tmp_ivl_8093;
  new_AGEMA_signal_3591 <= tmp_ivl_8100(1);
  n3733 <= tmp_ivl_8100(0);
  tmp_ivl_8100 <= LPM_d0_ivl_8104(0 + 1 downto 0);
  tmp_ivl_8106 <= state_in_s1(211);
  tmp_ivl_8108 <= state_in_s0(211);
  tmp_ivl_8109 <= tmp_ivl_8106 & tmp_ivl_8108;
  LPM_q_ivl_8112 <= tmp_ivl_8114 & tmp_ivl_8109;
  tmp_ivl_8117 <= z4(43);
  tmp_ivl_8118 <= new_AGEMA_signal_3148 & tmp_ivl_8117;
  LPM_q_ivl_8121 <= tmp_ivl_8123 & tmp_ivl_8118;
  new_AGEMA_signal_3302 <= tmp_ivl_8125(1);
  n3646 <= tmp_ivl_8125(0);
  tmp_ivl_8125 <= LPM_d0_ivl_8129(0 + 1 downto 0);
  tmp_ivl_8131 <= state_in_s1(275);
  tmp_ivl_8133 <= state_in_s0(275);
  tmp_ivl_8134 <= tmp_ivl_8131 & tmp_ivl_8133;
  LPM_q_ivl_8137 <= tmp_ivl_8139 & tmp_ivl_8134;
  tmp_ivl_8141 <= new_AGEMA_signal_3302 & n3646;
  LPM_q_ivl_8144 <= tmp_ivl_8146 & tmp_ivl_8141;
  new_AGEMA_signal_3592 <= tmp_ivl_8148(1);
  n3730 <= tmp_ivl_8148(0);
  tmp_ivl_8148 <= LPM_d0_ivl_8152(0 + 1 downto 0);
  tmp_ivl_8153 <= new_AGEMA_signal_3591 & n3733;
  LPM_q_ivl_8156 <= tmp_ivl_8158 & tmp_ivl_8153;
  tmp_ivl_8160 <= new_AGEMA_signal_3592 & n3730;
  LPM_q_ivl_8163 <= tmp_ivl_8165 & tmp_ivl_8160;
  new_AGEMA_signal_3893 <= tmp_ivl_8167(1);
  n3294 <= tmp_ivl_8167(0);
  tmp_ivl_8167 <= LPM_d0_ivl_8171(0 + 1 downto 0);
  tmp_ivl_8173 <= state_in_s1(250);
  tmp_ivl_8175 <= state_in_s0(250);
  tmp_ivl_8176 <= tmp_ivl_8173 & tmp_ivl_8175;
  LPM_q_ivl_8179 <= tmp_ivl_8181 & tmp_ivl_8176;
  tmp_ivl_8184 <= z4(2);
  tmp_ivl_8185 <= new_AGEMA_signal_3133 & tmp_ivl_8184;
  LPM_q_ivl_8188 <= tmp_ivl_8190 & tmp_ivl_8185;
  new_AGEMA_signal_3303 <= tmp_ivl_8192(1);
  n3706 <= tmp_ivl_8192(0);
  tmp_ivl_8192 <= LPM_d0_ivl_8196(0 + 1 downto 0);
  tmp_ivl_8198 <= state_in_s1(314);
  tmp_ivl_8200 <= state_in_s0(314);
  tmp_ivl_8201 <= tmp_ivl_8198 & tmp_ivl_8200;
  LPM_q_ivl_8204 <= tmp_ivl_8206 & tmp_ivl_8201;
  tmp_ivl_8208 <= new_AGEMA_signal_3303 & n3706;
  LPM_q_ivl_8211 <= tmp_ivl_8213 & tmp_ivl_8208;
  new_AGEMA_signal_3593 <= tmp_ivl_8215(1);
  n3360 <= tmp_ivl_8215(0);
  tmp_ivl_8215 <= LPM_d0_ivl_8219(0 + 1 downto 0);
  tmp_ivl_8220 <= new_AGEMA_signal_3893 & n3294;
  LPM_q_ivl_8223 <= tmp_ivl_8225 & tmp_ivl_8220;
  tmp_ivl_8227 <= new_AGEMA_signal_3593 & n3360;
  LPM_q_ivl_8230 <= tmp_ivl_8232 & tmp_ivl_8227;
  tmp_ivl_8234 <= tmp_ivl_8238(1);
  tmp_ivl_8236 <= tmp_ivl_8238(0);
  tmp_ivl_8238 <= LPM_d0_ivl_8242(0 + 1 downto 0);
  tmp_ivl_8244 <= state_in_s1(242);
  tmp_ivl_8246 <= state_in_s0(242);
  tmp_ivl_8247 <= tmp_ivl_8244 & tmp_ivl_8246;
  LPM_q_ivl_8250 <= tmp_ivl_8252 & tmp_ivl_8247;
  tmp_ivl_8255 <= z4(10);
  tmp_ivl_8256 <= new_AGEMA_signal_3112 & tmp_ivl_8255;
  LPM_q_ivl_8259 <= tmp_ivl_8261 & tmp_ivl_8256;
  new_AGEMA_signal_3304 <= tmp_ivl_8263(1);
  n3396 <= tmp_ivl_8263(0);
  tmp_ivl_8263 <= LPM_d0_ivl_8267(0 + 1 downto 0);
  tmp_ivl_8269 <= state_in_s1(306);
  tmp_ivl_8271 <= state_in_s0(306);
  tmp_ivl_8272 <= tmp_ivl_8269 & tmp_ivl_8271;
  LPM_q_ivl_8275 <= tmp_ivl_8277 & tmp_ivl_8272;
  tmp_ivl_8279 <= new_AGEMA_signal_3304 & n3396;
  LPM_q_ivl_8282 <= tmp_ivl_8284 & tmp_ivl_8279;
  new_AGEMA_signal_3594 <= tmp_ivl_8286(1);
  n3839 <= tmp_ivl_8286(0);
  tmp_ivl_8286 <= LPM_d0_ivl_8290(0 + 1 downto 0);
  tmp_ivl_8292 <= state_in_s1(212);
  tmp_ivl_8294 <= state_in_s0(212);
  tmp_ivl_8295 <= tmp_ivl_8292 & tmp_ivl_8294;
  LPM_q_ivl_8298 <= tmp_ivl_8300 & tmp_ivl_8295;
  tmp_ivl_8303 <= z4(44);
  tmp_ivl_8304 <= new_AGEMA_signal_3149 & tmp_ivl_8303;
  LPM_q_ivl_8307 <= tmp_ivl_8309 & tmp_ivl_8304;
  new_AGEMA_signal_3305 <= tmp_ivl_8311(1);
  n3692 <= tmp_ivl_8311(0);
  tmp_ivl_8311 <= LPM_d0_ivl_8315(0 + 1 downto 0);
  tmp_ivl_8317 <= state_in_s1(276);
  tmp_ivl_8319 <= state_in_s0(276);
  tmp_ivl_8320 <= tmp_ivl_8317 & tmp_ivl_8319;
  LPM_q_ivl_8323 <= tmp_ivl_8325 & tmp_ivl_8320;
  tmp_ivl_8327 <= new_AGEMA_signal_3305 & n3692;
  LPM_q_ivl_8330 <= tmp_ivl_8332 & tmp_ivl_8327;
  new_AGEMA_signal_3595 <= tmp_ivl_8334(1);
  n3836 <= tmp_ivl_8334(0);
  tmp_ivl_8334 <= LPM_d0_ivl_8338(0 + 1 downto 0);
  tmp_ivl_8339 <= new_AGEMA_signal_3594 & n3839;
  LPM_q_ivl_8342 <= tmp_ivl_8344 & tmp_ivl_8339;
  tmp_ivl_8346 <= new_AGEMA_signal_3595 & n3836;
  LPM_q_ivl_8349 <= tmp_ivl_8351 & tmp_ivl_8346;
  new_AGEMA_signal_3894 <= tmp_ivl_8353(1);
  n3295 <= tmp_ivl_8353(0);
  tmp_ivl_8353 <= LPM_d0_ivl_8357(0 + 1 downto 0);
  tmp_ivl_8359 <= state_in_s1(251);
  tmp_ivl_8361 <= state_in_s0(251);
  tmp_ivl_8362 <= tmp_ivl_8359 & tmp_ivl_8361;
  LPM_q_ivl_8365 <= tmp_ivl_8367 & tmp_ivl_8362;
  tmp_ivl_8370 <= z4(3);
  tmp_ivl_8371 <= new_AGEMA_signal_3144 & tmp_ivl_8370;
  LPM_q_ivl_8374 <= tmp_ivl_8376 & tmp_ivl_8371;
  new_AGEMA_signal_3306 <= tmp_ivl_8378(1);
  n3800 <= tmp_ivl_8378(0);
  tmp_ivl_8378 <= LPM_d0_ivl_8382(0 + 1 downto 0);
  tmp_ivl_8384 <= state_in_s1(315);
  tmp_ivl_8386 <= state_in_s0(315);
  tmp_ivl_8387 <= tmp_ivl_8384 & tmp_ivl_8386;
  LPM_q_ivl_8390 <= tmp_ivl_8392 & tmp_ivl_8387;
  tmp_ivl_8394 <= new_AGEMA_signal_3306 & n3800;
  LPM_q_ivl_8397 <= tmp_ivl_8399 & tmp_ivl_8394;
  new_AGEMA_signal_3596 <= tmp_ivl_8401(1);
  n3391 <= tmp_ivl_8401(0);
  tmp_ivl_8401 <= LPM_d0_ivl_8405(0 + 1 downto 0);
  tmp_ivl_8406 <= new_AGEMA_signal_3894 & n3295;
  LPM_q_ivl_8409 <= tmp_ivl_8411 & tmp_ivl_8406;
  tmp_ivl_8413 <= new_AGEMA_signal_3596 & n3391;
  LPM_q_ivl_8416 <= tmp_ivl_8418 & tmp_ivl_8413;
  tmp_ivl_8420 <= tmp_ivl_8424(1);
  tmp_ivl_8422 <= tmp_ivl_8424(0);
  tmp_ivl_8424 <= LPM_d0_ivl_8428(0 + 1 downto 0);
  tmp_ivl_8430 <= state_in_s1(243);
  tmp_ivl_8432 <= state_in_s0(243);
  tmp_ivl_8433 <= tmp_ivl_8430 & tmp_ivl_8432;
  LPM_q_ivl_8436 <= tmp_ivl_8438 & tmp_ivl_8433;
  tmp_ivl_8441 <= z4(11);
  tmp_ivl_8442 <= new_AGEMA_signal_3113 & tmp_ivl_8441;
  LPM_q_ivl_8445 <= tmp_ivl_8447 & tmp_ivl_8442;
  new_AGEMA_signal_3307 <= tmp_ivl_8449(1);
  n3438 <= tmp_ivl_8449(0);
  tmp_ivl_8449 <= LPM_d0_ivl_8453(0 + 1 downto 0);
  tmp_ivl_8455 <= state_in_s1(307);
  tmp_ivl_8457 <= state_in_s0(307);
  tmp_ivl_8458 <= tmp_ivl_8455 & tmp_ivl_8457;
  LPM_q_ivl_8461 <= tmp_ivl_8463 & tmp_ivl_8458;
  tmp_ivl_8465 <= new_AGEMA_signal_3307 & n3438;
  LPM_q_ivl_8468 <= tmp_ivl_8470 & tmp_ivl_8465;
  new_AGEMA_signal_3597 <= tmp_ivl_8472(1);
  n3929 <= tmp_ivl_8472(0);
  tmp_ivl_8472 <= LPM_d0_ivl_8476(0 + 1 downto 0);
  tmp_ivl_8478 <= state_in_s1(213);
  tmp_ivl_8480 <= state_in_s0(213);
  tmp_ivl_8481 <= tmp_ivl_8478 & tmp_ivl_8480;
  LPM_q_ivl_8484 <= tmp_ivl_8486 & tmp_ivl_8481;
  tmp_ivl_8489 <= z4(45);
  tmp_ivl_8490 <= new_AGEMA_signal_3150 & tmp_ivl_8489;
  LPM_q_ivl_8493 <= tmp_ivl_8495 & tmp_ivl_8490;
  new_AGEMA_signal_3308 <= tmp_ivl_8497(1);
  n3783 <= tmp_ivl_8497(0);
  tmp_ivl_8497 <= LPM_d0_ivl_8501(0 + 1 downto 0);
  tmp_ivl_8503 <= state_in_s1(277);
  tmp_ivl_8505 <= state_in_s0(277);
  tmp_ivl_8506 <= tmp_ivl_8503 & tmp_ivl_8505;
  LPM_q_ivl_8509 <= tmp_ivl_8511 & tmp_ivl_8506;
  tmp_ivl_8513 <= new_AGEMA_signal_3308 & n3783;
  LPM_q_ivl_8516 <= tmp_ivl_8518 & tmp_ivl_8513;
  new_AGEMA_signal_3598 <= tmp_ivl_8520(1);
  n3925 <= tmp_ivl_8520(0);
  tmp_ivl_8520 <= LPM_d0_ivl_8524(0 + 1 downto 0);
  tmp_ivl_8525 <= new_AGEMA_signal_3597 & n3929;
  LPM_q_ivl_8528 <= tmp_ivl_8530 & tmp_ivl_8525;
  tmp_ivl_8532 <= new_AGEMA_signal_3598 & n3925;
  LPM_q_ivl_8535 <= tmp_ivl_8537 & tmp_ivl_8532;
  new_AGEMA_signal_3895 <= tmp_ivl_8539(1);
  n3296 <= tmp_ivl_8539(0);
  tmp_ivl_8539 <= LPM_d0_ivl_8543(0 + 1 downto 0);
  tmp_ivl_8545 <= state_in_s1(252);
  tmp_ivl_8547 <= state_in_s0(252);
  tmp_ivl_8548 <= tmp_ivl_8545 & tmp_ivl_8547;
  LPM_q_ivl_8551 <= tmp_ivl_8553 & tmp_ivl_8548;
  tmp_ivl_8556 <= z4(4);
  tmp_ivl_8557 <= new_AGEMA_signal_3155 & tmp_ivl_8556;
  LPM_q_ivl_8560 <= tmp_ivl_8562 & tmp_ivl_8557;
  new_AGEMA_signal_3309 <= tmp_ivl_8564(1);
  n3888 <= tmp_ivl_8564(0);
  tmp_ivl_8564 <= LPM_d0_ivl_8568(0 + 1 downto 0);
  tmp_ivl_8570 <= state_in_s1(316);
  tmp_ivl_8572 <= state_in_s0(316);
  tmp_ivl_8573 <= tmp_ivl_8570 & tmp_ivl_8572;
  LPM_q_ivl_8576 <= tmp_ivl_8578 & tmp_ivl_8573;
  tmp_ivl_8580 <= new_AGEMA_signal_3309 & n3888;
  LPM_q_ivl_8583 <= tmp_ivl_8585 & tmp_ivl_8580;
  new_AGEMA_signal_3599 <= tmp_ivl_8587(1);
  n3454 <= tmp_ivl_8587(0);
  tmp_ivl_8587 <= LPM_d0_ivl_8591(0 + 1 downto 0);
  tmp_ivl_8592 <= new_AGEMA_signal_3895 & n3296;
  LPM_q_ivl_8595 <= tmp_ivl_8597 & tmp_ivl_8592;
  tmp_ivl_8599 <= new_AGEMA_signal_3599 & n3454;
  LPM_q_ivl_8602 <= tmp_ivl_8604 & tmp_ivl_8599;
  tmp_ivl_8606 <= tmp_ivl_8610(1);
  tmp_ivl_8608 <= tmp_ivl_8610(0);
  tmp_ivl_8610 <= LPM_d0_ivl_8614(0 + 1 downto 0);
  tmp_ivl_8616 <= state_in_s1(235);
  tmp_ivl_8618 <= state_in_s0(235);
  tmp_ivl_8619 <= tmp_ivl_8616 & tmp_ivl_8618;
  LPM_q_ivl_8622 <= tmp_ivl_8624 & tmp_ivl_8619;
  tmp_ivl_8627 <= z4(19);
  tmp_ivl_8628 <= new_AGEMA_signal_3121 & tmp_ivl_8627;
  LPM_q_ivl_8631 <= tmp_ivl_8633 & tmp_ivl_8628;
  new_AGEMA_signal_3310 <= tmp_ivl_8635(1);
  n3355 <= tmp_ivl_8635(0);
  tmp_ivl_8635 <= LPM_d0_ivl_8639(0 + 1 downto 0);
  tmp_ivl_8641 <= state_in_s1(299);
  tmp_ivl_8643 <= state_in_s0(299);
  tmp_ivl_8644 <= tmp_ivl_8641 & tmp_ivl_8643;
  LPM_q_ivl_8647 <= tmp_ivl_8649 & tmp_ivl_8644;
  tmp_ivl_8651 <= new_AGEMA_signal_3310 & n3355;
  LPM_q_ivl_8654 <= tmp_ivl_8656 & tmp_ivl_8651;
  new_AGEMA_signal_3600 <= tmp_ivl_8658(1);
  n3660 <= tmp_ivl_8658(0);
  tmp_ivl_8658 <= LPM_d0_ivl_8662(0 + 1 downto 0);
  tmp_ivl_8664 <= state_in_s1(205);
  tmp_ivl_8666 <= state_in_s0(205);
  tmp_ivl_8667 <= tmp_ivl_8664 & tmp_ivl_8666;
  LPM_q_ivl_8670 <= tmp_ivl_8672 & tmp_ivl_8667;
  tmp_ivl_8675 <= z4(53);
  tmp_ivl_8676 <= new_AGEMA_signal_3159 & tmp_ivl_8675;
  LPM_q_ivl_8679 <= tmp_ivl_8681 & tmp_ivl_8676;
  new_AGEMA_signal_3311 <= tmp_ivl_8683(1);
  n3566 <= tmp_ivl_8683(0);
  tmp_ivl_8683 <= LPM_d0_ivl_8687(0 + 1 downto 0);
  tmp_ivl_8689 <= state_in_s1(269);
  tmp_ivl_8691 <= state_in_s0(269);
  tmp_ivl_8692 <= tmp_ivl_8689 & tmp_ivl_8691;
  LPM_q_ivl_8695 <= tmp_ivl_8697 & tmp_ivl_8692;
  tmp_ivl_8699 <= new_AGEMA_signal_3311 & n3566;
  LPM_q_ivl_8702 <= tmp_ivl_8704 & tmp_ivl_8699;
  new_AGEMA_signal_3601 <= tmp_ivl_8706(1);
  n3625 <= tmp_ivl_8706(0);
  tmp_ivl_8706 <= LPM_d0_ivl_8710(0 + 1 downto 0);
  tmp_ivl_8711 <= new_AGEMA_signal_3600 & n3660;
  LPM_q_ivl_8714 <= tmp_ivl_8716 & tmp_ivl_8711;
  tmp_ivl_8718 <= new_AGEMA_signal_3601 & n3625;
  LPM_q_ivl_8721 <= tmp_ivl_8723 & tmp_ivl_8718;
  new_AGEMA_signal_3896 <= tmp_ivl_8725(1);
  n3297 <= tmp_ivl_8725(0);
  tmp_ivl_8725 <= LPM_d0_ivl_8729(0 + 1 downto 0);
  tmp_ivl_8731 <= state_in_s1(244);
  tmp_ivl_8733 <= state_in_s0(244);
  tmp_ivl_8734 <= tmp_ivl_8731 & tmp_ivl_8733;
  LPM_q_ivl_8737 <= tmp_ivl_8739 & tmp_ivl_8734;
  tmp_ivl_8742 <= z4(12);
  tmp_ivl_8743 <= new_AGEMA_signal_3114 & tmp_ivl_8742;
  LPM_q_ivl_8746 <= tmp_ivl_8748 & tmp_ivl_8743;
  new_AGEMA_signal_3312 <= tmp_ivl_8750(1);
  n3493 <= tmp_ivl_8750(0);
  tmp_ivl_8750 <= LPM_d0_ivl_8754(0 + 1 downto 0);
  tmp_ivl_8756 <= state_in_s1(308);
  tmp_ivl_8758 <= state_in_s0(308);
  tmp_ivl_8759 <= tmp_ivl_8756 & tmp_ivl_8758;
  LPM_q_ivl_8762 <= tmp_ivl_8764 & tmp_ivl_8759;
  tmp_ivl_8766 <= new_AGEMA_signal_3312 & n3493;
  LPM_q_ivl_8769 <= tmp_ivl_8771 & tmp_ivl_8766;
  new_AGEMA_signal_3602 <= tmp_ivl_8773(1);
  n3304 <= tmp_ivl_8773(0);
  tmp_ivl_8773 <= LPM_d0_ivl_8777(0 + 1 downto 0);
  tmp_ivl_8778 <= new_AGEMA_signal_3896 & n3297;
  LPM_q_ivl_8781 <= tmp_ivl_8783 & tmp_ivl_8778;
  tmp_ivl_8785 <= new_AGEMA_signal_3602 & n3304;
  LPM_q_ivl_8788 <= tmp_ivl_8790 & tmp_ivl_8785;
  tmp_ivl_8792 <= tmp_ivl_8796(1);
  tmp_ivl_8794 <= tmp_ivl_8796(0);
  tmp_ivl_8796 <= LPM_d0_ivl_8800(0 + 1 downto 0);
  tmp_ivl_8802 <= state_in_s1(214);
  tmp_ivl_8804 <= state_in_s0(214);
  tmp_ivl_8805 <= tmp_ivl_8802 & tmp_ivl_8804;
  LPM_q_ivl_8808 <= tmp_ivl_8810 & tmp_ivl_8805;
  tmp_ivl_8813 <= z4(46);
  tmp_ivl_8814 <= new_AGEMA_signal_3151 & tmp_ivl_8813;
  LPM_q_ivl_8817 <= tmp_ivl_8819 & tmp_ivl_8814;
  new_AGEMA_signal_3313 <= tmp_ivl_8821(1);
  n3844 <= tmp_ivl_8821(0);
  tmp_ivl_8821 <= LPM_d0_ivl_8825(0 + 1 downto 0);
  tmp_ivl_8827 <= state_in_s1(278);
  tmp_ivl_8829 <= state_in_s0(278);
  tmp_ivl_8830 <= tmp_ivl_8827 & tmp_ivl_8829;
  LPM_q_ivl_8833 <= tmp_ivl_8835 & tmp_ivl_8830;
  tmp_ivl_8837 <= new_AGEMA_signal_3313 & n3844;
  LPM_q_ivl_8840 <= tmp_ivl_8842 & tmp_ivl_8837;
  new_AGEMA_signal_3603 <= tmp_ivl_8844(1);
  n3687 <= tmp_ivl_8844(0);
  tmp_ivl_8844 <= LPM_d0_ivl_8848(0 + 1 downto 0);
  tmp_ivl_8849 <= new_AGEMA_signal_3602 & n3304;
  LPM_q_ivl_8852 <= tmp_ivl_8854 & tmp_ivl_8849;
  tmp_ivl_8856 <= new_AGEMA_signal_3603 & n3687;
  LPM_q_ivl_8859 <= tmp_ivl_8861 & tmp_ivl_8856;
  new_AGEMA_signal_3897 <= tmp_ivl_8863(1);
  n3298 <= tmp_ivl_8863(0);
  tmp_ivl_8863 <= LPM_d0_ivl_8867(0 + 1 downto 0);
  tmp_ivl_8869 <= state_in_s1(253);
  tmp_ivl_8871 <= state_in_s0(253);
  tmp_ivl_8872 <= tmp_ivl_8869 & tmp_ivl_8871;
  LPM_q_ivl_8875 <= tmp_ivl_8877 & tmp_ivl_8872;
  tmp_ivl_8880 <= z4(5);
  tmp_ivl_8881 <= new_AGEMA_signal_3166 & tmp_ivl_8880;
  LPM_q_ivl_8884 <= tmp_ivl_8886 & tmp_ivl_8881;
  new_AGEMA_signal_3314 <= tmp_ivl_8888(1);
  n3738 <= tmp_ivl_8888(0);
  tmp_ivl_8888 <= LPM_d0_ivl_8892(0 + 1 downto 0);
  tmp_ivl_8894 <= state_in_s1(317);
  tmp_ivl_8896 <= state_in_s0(317);
  tmp_ivl_8897 <= tmp_ivl_8894 & tmp_ivl_8896;
  LPM_q_ivl_8900 <= tmp_ivl_8902 & tmp_ivl_8897;
  tmp_ivl_8904 <= new_AGEMA_signal_3314 & n3738;
  LPM_q_ivl_8907 <= tmp_ivl_8909 & tmp_ivl_8904;
  new_AGEMA_signal_3604 <= tmp_ivl_8911(1);
  n3508 <= tmp_ivl_8911(0);
  tmp_ivl_8911 <= LPM_d0_ivl_8915(0 + 1 downto 0);
  tmp_ivl_8916 <= new_AGEMA_signal_3897 & n3298;
  LPM_q_ivl_8919 <= tmp_ivl_8921 & tmp_ivl_8916;
  tmp_ivl_8923 <= new_AGEMA_signal_3604 & n3508;
  LPM_q_ivl_8926 <= tmp_ivl_8928 & tmp_ivl_8923;
  tmp_ivl_8930 <= tmp_ivl_8934(1);
  tmp_ivl_8932 <= tmp_ivl_8934(0);
  tmp_ivl_8934 <= LPM_d0_ivl_8938(0 + 1 downto 0);
  tmp_ivl_8940 <= state_in_s1(236);
  tmp_ivl_8942 <= state_in_s0(236);
  tmp_ivl_8943 <= tmp_ivl_8940 & tmp_ivl_8942;
  LPM_q_ivl_8946 <= tmp_ivl_8948 & tmp_ivl_8943;
  tmp_ivl_8951 <= z4(20);
  tmp_ivl_8952 <= new_AGEMA_signal_3123 & tmp_ivl_8951;
  LPM_q_ivl_8955 <= tmp_ivl_8957 & tmp_ivl_8952;
  new_AGEMA_signal_3315 <= tmp_ivl_8959(1);
  n3439 <= tmp_ivl_8959(0);
  tmp_ivl_8959 <= LPM_d0_ivl_8963(0 + 1 downto 0);
  tmp_ivl_8965 <= state_in_s1(300);
  tmp_ivl_8967 <= state_in_s0(300);
  tmp_ivl_8968 <= tmp_ivl_8965 & tmp_ivl_8967;
  LPM_q_ivl_8971 <= tmp_ivl_8973 & tmp_ivl_8968;
  tmp_ivl_8975 <= new_AGEMA_signal_3315 & n3439;
  LPM_q_ivl_8978 <= tmp_ivl_8980 & tmp_ivl_8975;
  new_AGEMA_signal_3605 <= tmp_ivl_8982(1);
  n3729 <= tmp_ivl_8982(0);
  tmp_ivl_8982 <= LPM_d0_ivl_8986(0 + 1 downto 0);
  tmp_ivl_8988 <= state_in_s1(206);
  tmp_ivl_8990 <= state_in_s0(206);
  tmp_ivl_8991 <= tmp_ivl_8988 & tmp_ivl_8990;
  LPM_q_ivl_8994 <= tmp_ivl_8996 & tmp_ivl_8991;
  tmp_ivl_8999 <= z4(54);
  tmp_ivl_9000 <= new_AGEMA_signal_3160 & tmp_ivl_8999;
  LPM_q_ivl_9003 <= tmp_ivl_9005 & tmp_ivl_9000;
  new_AGEMA_signal_3316 <= tmp_ivl_9007(1);
  n3582 <= tmp_ivl_9007(0);
  tmp_ivl_9007 <= LPM_d0_ivl_9011(0 + 1 downto 0);
  tmp_ivl_9013 <= state_in_s1(270);
  tmp_ivl_9015 <= state_in_s0(270);
  tmp_ivl_9016 <= tmp_ivl_9013 & tmp_ivl_9015;
  LPM_q_ivl_9019 <= tmp_ivl_9021 & tmp_ivl_9016;
  tmp_ivl_9023 <= new_AGEMA_signal_3316 & n3582;
  LPM_q_ivl_9026 <= tmp_ivl_9028 & tmp_ivl_9023;
  new_AGEMA_signal_3606 <= tmp_ivl_9030(1);
  n3457 <= tmp_ivl_9030(0);
  tmp_ivl_9030 <= LPM_d0_ivl_9034(0 + 1 downto 0);
  tmp_ivl_9035 <= new_AGEMA_signal_3605 & n3729;
  LPM_q_ivl_9038 <= tmp_ivl_9040 & tmp_ivl_9035;
  tmp_ivl_9042 <= new_AGEMA_signal_3606 & n3457;
  LPM_q_ivl_9045 <= tmp_ivl_9047 & tmp_ivl_9042;
  new_AGEMA_signal_3898 <= tmp_ivl_9049(1);
  n3299 <= tmp_ivl_9049(0);
  tmp_ivl_9049 <= LPM_d0_ivl_9053(0 + 1 downto 0);
  tmp_ivl_9055 <= state_in_s1(245);
  tmp_ivl_9057 <= state_in_s0(245);
  tmp_ivl_9058 <= tmp_ivl_9055 & tmp_ivl_9057;
  LPM_q_ivl_9061 <= tmp_ivl_9063 & tmp_ivl_9058;
  tmp_ivl_9066 <= z4(13);
  tmp_ivl_9067 <= new_AGEMA_signal_3115 & tmp_ivl_9066;
  LPM_q_ivl_9070 <= tmp_ivl_9072 & tmp_ivl_9067;
  new_AGEMA_signal_3317 <= tmp_ivl_9074(1);
  n3404 <= tmp_ivl_9074(0);
  tmp_ivl_9074 <= LPM_d0_ivl_9078(0 + 1 downto 0);
  tmp_ivl_9080 <= state_in_s1(309);
  tmp_ivl_9082 <= state_in_s0(309);
  tmp_ivl_9083 <= tmp_ivl_9080 & tmp_ivl_9082;
  LPM_q_ivl_9086 <= tmp_ivl_9088 & tmp_ivl_9083;
  tmp_ivl_9090 <= new_AGEMA_signal_3317 & n3404;
  LPM_q_ivl_9093 <= tmp_ivl_9095 & tmp_ivl_9090;
  new_AGEMA_signal_3607 <= tmp_ivl_9097(1);
  n3306 <= tmp_ivl_9097(0);
  tmp_ivl_9097 <= LPM_d0_ivl_9101(0 + 1 downto 0);
  tmp_ivl_9102 <= new_AGEMA_signal_3898 & n3299;
  LPM_q_ivl_9105 <= tmp_ivl_9107 & tmp_ivl_9102;
  tmp_ivl_9109 <= new_AGEMA_signal_3607 & n3306;
  LPM_q_ivl_9112 <= tmp_ivl_9114 & tmp_ivl_9109;
  tmp_ivl_9116 <= tmp_ivl_9120(1);
  tmp_ivl_9118 <= tmp_ivl_9120(0);
  tmp_ivl_9120 <= LPM_d0_ivl_9124(0 + 1 downto 0);
  tmp_ivl_9126 <= state_in_s1(215);
  tmp_ivl_9128 <= state_in_s0(215);
  tmp_ivl_9129 <= tmp_ivl_9126 & tmp_ivl_9128;
  LPM_q_ivl_9132 <= tmp_ivl_9134 & tmp_ivl_9129;
  tmp_ivl_9137 <= z4(47);
  tmp_ivl_9138 <= new_AGEMA_signal_3152 & tmp_ivl_9137;
  LPM_q_ivl_9141 <= tmp_ivl_9143 & tmp_ivl_9138;
  new_AGEMA_signal_3318 <= tmp_ivl_9145(1);
  n3354 <= tmp_ivl_9145(0);
  tmp_ivl_9145 <= LPM_d0_ivl_9149(0 + 1 downto 0);
  tmp_ivl_9151 <= state_in_s1(279);
  tmp_ivl_9153 <= state_in_s0(279);
  tmp_ivl_9154 <= tmp_ivl_9151 & tmp_ivl_9153;
  LPM_q_ivl_9157 <= tmp_ivl_9159 & tmp_ivl_9154;
  tmp_ivl_9161 <= new_AGEMA_signal_3318 & n3354;
  LPM_q_ivl_9164 <= tmp_ivl_9166 & tmp_ivl_9161;
  new_AGEMA_signal_3608 <= tmp_ivl_9168(1);
  n3777 <= tmp_ivl_9168(0);
  tmp_ivl_9168 <= LPM_d0_ivl_9172(0 + 1 downto 0);
  tmp_ivl_9173 <= new_AGEMA_signal_3607 & n3306;
  LPM_q_ivl_9176 <= tmp_ivl_9178 & tmp_ivl_9173;
  tmp_ivl_9180 <= new_AGEMA_signal_3608 & n3777;
  LPM_q_ivl_9183 <= tmp_ivl_9185 & tmp_ivl_9180;
  new_AGEMA_signal_3899 <= tmp_ivl_9187(1);
  n3300 <= tmp_ivl_9187(0);
  tmp_ivl_9187 <= LPM_d0_ivl_9191(0 + 1 downto 0);
  tmp_ivl_9193 <= state_in_s1(254);
  tmp_ivl_9195 <= state_in_s0(254);
  tmp_ivl_9196 <= tmp_ivl_9193 & tmp_ivl_9195;
  LPM_q_ivl_9199 <= tmp_ivl_9201 & tmp_ivl_9196;
  tmp_ivl_9204 <= z4(6);
  tmp_ivl_9205 <= new_AGEMA_signal_3171 & tmp_ivl_9204;
  LPM_q_ivl_9208 <= tmp_ivl_9210 & tmp_ivl_9205;
  new_AGEMA_signal_3319 <= tmp_ivl_9212(1);
  n3757 <= tmp_ivl_9212(0);
  tmp_ivl_9212 <= LPM_d0_ivl_9216(0 + 1 downto 0);
  tmp_ivl_9218 <= state_in_s1(318);
  tmp_ivl_9220 <= state_in_s0(318);
  tmp_ivl_9221 <= tmp_ivl_9218 & tmp_ivl_9220;
  LPM_q_ivl_9224 <= tmp_ivl_9226 & tmp_ivl_9221;
  tmp_ivl_9228 <= new_AGEMA_signal_3319 & n3757;
  LPM_q_ivl_9231 <= tmp_ivl_9233 & tmp_ivl_9228;
  new_AGEMA_signal_3609 <= tmp_ivl_9235(1);
  n3561 <= tmp_ivl_9235(0);
  tmp_ivl_9235 <= LPM_d0_ivl_9239(0 + 1 downto 0);
  tmp_ivl_9240 <= new_AGEMA_signal_3899 & n3300;
  LPM_q_ivl_9243 <= tmp_ivl_9245 & tmp_ivl_9240;
  tmp_ivl_9247 <= new_AGEMA_signal_3609 & n3561;
  LPM_q_ivl_9250 <= tmp_ivl_9252 & tmp_ivl_9247;
  tmp_ivl_9254 <= tmp_ivl_9258(1);
  tmp_ivl_9256 <= tmp_ivl_9258(0);
  tmp_ivl_9258 <= LPM_d0_ivl_9262(0 + 1 downto 0);
  tmp_ivl_9264 <= state_in_s1(223);
  tmp_ivl_9266 <= state_in_s0(223);
  tmp_ivl_9267 <= tmp_ivl_9264 & tmp_ivl_9266;
  LPM_q_ivl_9270 <= tmp_ivl_9272 & tmp_ivl_9267;
  tmp_ivl_9275 <= z4(39);
  tmp_ivl_9276 <= new_AGEMA_signal_3143 & tmp_ivl_9275;
  LPM_q_ivl_9279 <= tmp_ivl_9281 & tmp_ivl_9276;
  new_AGEMA_signal_3320 <= tmp_ivl_9283(1);
  n3526 <= tmp_ivl_9283(0);
  tmp_ivl_9283 <= LPM_d0_ivl_9287(0 + 1 downto 0);
  tmp_ivl_9289 <= state_in_s1(287);
  tmp_ivl_9291 <= state_in_s0(287);
  tmp_ivl_9292 <= tmp_ivl_9289 & tmp_ivl_9291;
  LPM_q_ivl_9295 <= tmp_ivl_9297 & tmp_ivl_9292;
  tmp_ivl_9299 <= new_AGEMA_signal_3320 & n3526;
  LPM_q_ivl_9302 <= tmp_ivl_9304 & tmp_ivl_9299;
  new_AGEMA_signal_3610 <= tmp_ivl_9306(1);
  n3686 <= tmp_ivl_9306(0);
  tmp_ivl_9306 <= LPM_d0_ivl_9310(0 + 1 downto 0);
  tmp_ivl_9311 <= new_AGEMA_signal_3591 & n3733;
  LPM_q_ivl_9314 <= tmp_ivl_9316 & tmp_ivl_9311;
  tmp_ivl_9318 <= new_AGEMA_signal_3610 & n3686;
  LPM_q_ivl_9321 <= tmp_ivl_9323 & tmp_ivl_9318;
  new_AGEMA_signal_3900 <= tmp_ivl_9325(1);
  n3301 <= tmp_ivl_9325(0);
  tmp_ivl_9325 <= LPM_d0_ivl_9329(0 + 1 downto 0);
  tmp_ivl_9331 <= state_in_s1(216);
  tmp_ivl_9333 <= state_in_s0(216);
  tmp_ivl_9334 <= tmp_ivl_9331 & tmp_ivl_9333;
  LPM_q_ivl_9337 <= tmp_ivl_9339 & tmp_ivl_9334;
  tmp_ivl_9342 <= z4(32);
  tmp_ivl_9343 <= new_AGEMA_signal_3136 & tmp_ivl_9342;
  LPM_q_ivl_9346 <= tmp_ivl_9348 & tmp_ivl_9343;
  new_AGEMA_signal_3321 <= tmp_ivl_9350(1);
  n3603 <= tmp_ivl_9350(0);
  tmp_ivl_9350 <= LPM_d0_ivl_9354(0 + 1 downto 0);
  tmp_ivl_9356 <= state_in_s1(280);
  tmp_ivl_9358 <= state_in_s0(280);
  tmp_ivl_9359 <= tmp_ivl_9356 & tmp_ivl_9358;
  LPM_q_ivl_9362 <= tmp_ivl_9364 & tmp_ivl_9359;
  tmp_ivl_9366 <= new_AGEMA_signal_3321 & n3603;
  LPM_q_ivl_9369 <= tmp_ivl_9371 & tmp_ivl_9366;
  new_AGEMA_signal_3611 <= tmp_ivl_9373(1);
  n3511 <= tmp_ivl_9373(0);
  tmp_ivl_9373 <= LPM_d0_ivl_9377(0 + 1 downto 0);
  tmp_ivl_9378 <= new_AGEMA_signal_3900 & n3301;
  LPM_q_ivl_9381 <= tmp_ivl_9383 & tmp_ivl_9378;
  tmp_ivl_9385 <= new_AGEMA_signal_3611 & n3511;
  LPM_q_ivl_9388 <= tmp_ivl_9390 & tmp_ivl_9385;
  tmp_ivl_9392 <= tmp_ivl_9396(1);
  tmp_ivl_9394 <= tmp_ivl_9396(0);
  tmp_ivl_9396 <= LPM_d0_ivl_9400(0 + 1 downto 0);
  tmp_ivl_9402 <= state_in_s1(208);
  tmp_ivl_9404 <= state_in_s0(208);
  tmp_ivl_9405 <= tmp_ivl_9402 & tmp_ivl_9404;
  LPM_q_ivl_9408 <= tmp_ivl_9410 & tmp_ivl_9405;
  tmp_ivl_9413 <= z4(40);
  tmp_ivl_9414 <= new_AGEMA_signal_3145 & tmp_ivl_9413;
  LPM_q_ivl_9417 <= tmp_ivl_9419 & tmp_ivl_9414;
  new_AGEMA_signal_3322 <= tmp_ivl_9421(1);
  n3550 <= tmp_ivl_9421(0);
  tmp_ivl_9421 <= LPM_d0_ivl_9425(0 + 1 downto 0);
  tmp_ivl_9427 <= state_in_s1(272);
  tmp_ivl_9429 <= state_in_s0(272);
  tmp_ivl_9430 <= tmp_ivl_9427 & tmp_ivl_9429;
  LPM_q_ivl_9433 <= tmp_ivl_9435 & tmp_ivl_9430;
  tmp_ivl_9437 <= new_AGEMA_signal_3322 & n3550;
  LPM_q_ivl_9440 <= tmp_ivl_9442 & tmp_ivl_9437;
  new_AGEMA_signal_3612 <= tmp_ivl_9444(1);
  n3776 <= tmp_ivl_9444(0);
  tmp_ivl_9444 <= LPM_d0_ivl_9448(0 + 1 downto 0);
  tmp_ivl_9449 <= new_AGEMA_signal_3594 & n3839;
  LPM_q_ivl_9452 <= tmp_ivl_9454 & tmp_ivl_9449;
  tmp_ivl_9456 <= new_AGEMA_signal_3612 & n3776;
  LPM_q_ivl_9459 <= tmp_ivl_9461 & tmp_ivl_9456;
  new_AGEMA_signal_3901 <= tmp_ivl_9463(1);
  n3302 <= tmp_ivl_9463(0);
  tmp_ivl_9463 <= LPM_d0_ivl_9467(0 + 1 downto 0);
  tmp_ivl_9469 <= state_in_s1(217);
  tmp_ivl_9471 <= state_in_s0(217);
  tmp_ivl_9472 <= tmp_ivl_9469 & tmp_ivl_9471;
  LPM_q_ivl_9475 <= tmp_ivl_9477 & tmp_ivl_9472;
  tmp_ivl_9480 <= z4(33);
  tmp_ivl_9481 <= new_AGEMA_signal_3137 & tmp_ivl_9480;
  LPM_q_ivl_9484 <= tmp_ivl_9486 & tmp_ivl_9481;
  new_AGEMA_signal_3323 <= tmp_ivl_9488(1);
  n3613 <= tmp_ivl_9488(0);
  tmp_ivl_9488 <= LPM_d0_ivl_9492(0 + 1 downto 0);
  tmp_ivl_9494 <= state_in_s1(281);
  tmp_ivl_9496 <= state_in_s0(281);
  tmp_ivl_9497 <= tmp_ivl_9494 & tmp_ivl_9496;
  LPM_q_ivl_9500 <= tmp_ivl_9502 & tmp_ivl_9497;
  tmp_ivl_9504 <= new_AGEMA_signal_3323 & n3613;
  LPM_q_ivl_9507 <= tmp_ivl_9509 & tmp_ivl_9504;
  new_AGEMA_signal_3613 <= tmp_ivl_9511(1);
  n3559 <= tmp_ivl_9511(0);
  tmp_ivl_9511 <= LPM_d0_ivl_9515(0 + 1 downto 0);
  tmp_ivl_9516 <= new_AGEMA_signal_3901 & n3302;
  LPM_q_ivl_9519 <= tmp_ivl_9521 & tmp_ivl_9516;
  tmp_ivl_9523 <= new_AGEMA_signal_3613 & n3559;
  LPM_q_ivl_9526 <= tmp_ivl_9528 & tmp_ivl_9523;
  tmp_ivl_9530 <= tmp_ivl_9534(1);
  tmp_ivl_9532 <= tmp_ivl_9534(0);
  tmp_ivl_9534 <= LPM_d0_ivl_9538(0 + 1 downto 0);
  tmp_ivl_9540 <= state_in_s1(209);
  tmp_ivl_9542 <= state_in_s0(209);
  tmp_ivl_9543 <= tmp_ivl_9540 & tmp_ivl_9542;
  LPM_q_ivl_9546 <= tmp_ivl_9548 & tmp_ivl_9543;
  tmp_ivl_9551 <= z4(41);
  tmp_ivl_9552 <= new_AGEMA_signal_3146 & tmp_ivl_9551;
  LPM_q_ivl_9555 <= tmp_ivl_9557 & tmp_ivl_9552;
  new_AGEMA_signal_3324 <= tmp_ivl_9559(1);
  n3605 <= tmp_ivl_9559(0);
  tmp_ivl_9559 <= LPM_d0_ivl_9563(0 + 1 downto 0);
  tmp_ivl_9565 <= state_in_s1(273);
  tmp_ivl_9567 <= state_in_s0(273);
  tmp_ivl_9568 <= tmp_ivl_9565 & tmp_ivl_9567;
  LPM_q_ivl_9571 <= tmp_ivl_9573 & tmp_ivl_9568;
  tmp_ivl_9575 <= new_AGEMA_signal_3324 & n3605;
  LPM_q_ivl_9578 <= tmp_ivl_9580 & tmp_ivl_9575;
  new_AGEMA_signal_3614 <= tmp_ivl_9582(1);
  n3867 <= tmp_ivl_9582(0);
  tmp_ivl_9582 <= LPM_d0_ivl_9586(0 + 1 downto 0);
  tmp_ivl_9587 <= new_AGEMA_signal_3597 & n3929;
  LPM_q_ivl_9590 <= tmp_ivl_9592 & tmp_ivl_9587;
  tmp_ivl_9594 <= new_AGEMA_signal_3614 & n3867;
  LPM_q_ivl_9597 <= tmp_ivl_9599 & tmp_ivl_9594;
  new_AGEMA_signal_3902 <= tmp_ivl_9601(1);
  n3303 <= tmp_ivl_9601(0);
  tmp_ivl_9601 <= LPM_d0_ivl_9605(0 + 1 downto 0);
  tmp_ivl_9607 <= state_in_s1(218);
  tmp_ivl_9609 <= state_in_s0(218);
  tmp_ivl_9610 <= tmp_ivl_9607 & tmp_ivl_9609;
  LPM_q_ivl_9613 <= tmp_ivl_9615 & tmp_ivl_9610;
  tmp_ivl_9618 <= z4(34);
  tmp_ivl_9619 <= new_AGEMA_signal_3138 & tmp_ivl_9618;
  LPM_q_ivl_9622 <= tmp_ivl_9624 & tmp_ivl_9619;
  new_AGEMA_signal_3325 <= tmp_ivl_9626(1);
  n3568 <= tmp_ivl_9626(0);
  tmp_ivl_9626 <= LPM_d0_ivl_9630(0 + 1 downto 0);
  tmp_ivl_9632 <= state_in_s1(282);
  tmp_ivl_9634 <= state_in_s0(282);
  tmp_ivl_9635 <= tmp_ivl_9632 & tmp_ivl_9634;
  LPM_q_ivl_9638 <= tmp_ivl_9640 & tmp_ivl_9635;
  tmp_ivl_9642 <= new_AGEMA_signal_3325 & n3568;
  LPM_q_ivl_9645 <= tmp_ivl_9647 & tmp_ivl_9642;
  new_AGEMA_signal_3615 <= tmp_ivl_9649(1);
  n3422 <= tmp_ivl_9649(0);
  tmp_ivl_9649 <= LPM_d0_ivl_9653(0 + 1 downto 0);
  tmp_ivl_9654 <= new_AGEMA_signal_3902 & n3303;
  LPM_q_ivl_9657 <= tmp_ivl_9659 & tmp_ivl_9654;
  tmp_ivl_9661 <= new_AGEMA_signal_3615 & n3422;
  LPM_q_ivl_9664 <= tmp_ivl_9666 & tmp_ivl_9661;
  tmp_ivl_9668 <= tmp_ivl_9672(1);
  tmp_ivl_9670 <= tmp_ivl_9672(0);
  tmp_ivl_9672 <= LPM_d0_ivl_9676(0 + 1 downto 0);
  tmp_ivl_9677 <= new_AGEMA_signal_3589 & n3661;
  LPM_q_ivl_9680 <= tmp_ivl_9682 & tmp_ivl_9677;
  tmp_ivl_9684 <= new_AGEMA_signal_3602 & n3304;
  LPM_q_ivl_9687 <= tmp_ivl_9689 & tmp_ivl_9684;
  new_AGEMA_signal_3903 <= tmp_ivl_9691(1);
  n3305 <= tmp_ivl_9691(0);
  tmp_ivl_9691 <= LPM_d0_ivl_9695(0 + 1 downto 0);
  tmp_ivl_9697 <= state_in_s1(219);
  tmp_ivl_9699 <= state_in_s0(219);
  tmp_ivl_9700 <= tmp_ivl_9697 & tmp_ivl_9699;
  LPM_q_ivl_9703 <= tmp_ivl_9705 & tmp_ivl_9700;
  tmp_ivl_9708 <= z4(35);
  tmp_ivl_9709 <= new_AGEMA_signal_3139 & tmp_ivl_9708;
  LPM_q_ivl_9712 <= tmp_ivl_9714 & tmp_ivl_9709;
  new_AGEMA_signal_3326 <= tmp_ivl_9716(1);
  n3580 <= tmp_ivl_9716(0);
  tmp_ivl_9716 <= LPM_d0_ivl_9720(0 + 1 downto 0);
  tmp_ivl_9722 <= state_in_s1(283);
  tmp_ivl_9724 <= state_in_s0(283);
  tmp_ivl_9725 <= tmp_ivl_9722 & tmp_ivl_9724;
  LPM_q_ivl_9728 <= tmp_ivl_9730 & tmp_ivl_9725;
  tmp_ivl_9732 <= new_AGEMA_signal_3326 & n3580;
  LPM_q_ivl_9735 <= tmp_ivl_9737 & tmp_ivl_9732;
  new_AGEMA_signal_3616 <= tmp_ivl_9739(1);
  n3481 <= tmp_ivl_9739(0);
  tmp_ivl_9739 <= LPM_d0_ivl_9743(0 + 1 downto 0);
  tmp_ivl_9744 <= new_AGEMA_signal_3903 & n3305;
  LPM_q_ivl_9747 <= tmp_ivl_9749 & tmp_ivl_9744;
  tmp_ivl_9751 <= new_AGEMA_signal_3616 & n3481;
  LPM_q_ivl_9754 <= tmp_ivl_9756 & tmp_ivl_9751;
  tmp_ivl_9758 <= tmp_ivl_9762(1);
  tmp_ivl_9760 <= tmp_ivl_9762(0);
  tmp_ivl_9762 <= LPM_d0_ivl_9766(0 + 1 downto 0);
  tmp_ivl_9767 <= new_AGEMA_signal_3592 & n3730;
  LPM_q_ivl_9770 <= tmp_ivl_9772 & tmp_ivl_9767;
  tmp_ivl_9774 <= new_AGEMA_signal_3607 & n3306;
  LPM_q_ivl_9777 <= tmp_ivl_9779 & tmp_ivl_9774;
  new_AGEMA_signal_3904 <= tmp_ivl_9781(1);
  n3307 <= tmp_ivl_9781(0);
  tmp_ivl_9781 <= LPM_d0_ivl_9785(0 + 1 downto 0);
  tmp_ivl_9787 <= state_in_s1(220);
  tmp_ivl_9789 <= state_in_s0(220);
  tmp_ivl_9790 <= tmp_ivl_9787 & tmp_ivl_9789;
  LPM_q_ivl_9793 <= tmp_ivl_9795 & tmp_ivl_9790;
  tmp_ivl_9798 <= z4(36);
  tmp_ivl_9799 <= new_AGEMA_signal_3140 & tmp_ivl_9798;
  LPM_q_ivl_9802 <= tmp_ivl_9804 & tmp_ivl_9799;
  new_AGEMA_signal_3327 <= tmp_ivl_9806(1);
  n3418 <= tmp_ivl_9806(0);
  tmp_ivl_9806 <= LPM_d0_ivl_9810(0 + 1 downto 0);
  tmp_ivl_9812 <= state_in_s1(284);
  tmp_ivl_9814 <= state_in_s0(284);
  tmp_ivl_9815 <= tmp_ivl_9812 & tmp_ivl_9814;
  LPM_q_ivl_9818 <= tmp_ivl_9820 & tmp_ivl_9815;
  tmp_ivl_9822 <= new_AGEMA_signal_3327 & n3418;
  LPM_q_ivl_9825 <= tmp_ivl_9827 & tmp_ivl_9822;
  new_AGEMA_signal_3617 <= tmp_ivl_9829(1);
  n3538 <= tmp_ivl_9829(0);
  tmp_ivl_9829 <= LPM_d0_ivl_9833(0 + 1 downto 0);
  tmp_ivl_9834 <= new_AGEMA_signal_3904 & n3307;
  LPM_q_ivl_9837 <= tmp_ivl_9839 & tmp_ivl_9834;
  tmp_ivl_9841 <= new_AGEMA_signal_3617 & n3538;
  LPM_q_ivl_9844 <= tmp_ivl_9846 & tmp_ivl_9841;
  tmp_ivl_9848 <= tmp_ivl_9852(1);
  tmp_ivl_9850 <= tmp_ivl_9852(0);
  tmp_ivl_9852 <= LPM_d0_ivl_9856(0 + 1 downto 0);
  tmp_ivl_9858 <= state_in_s1(221);
  tmp_ivl_9860 <= state_in_s0(221);
  tmp_ivl_9861 <= tmp_ivl_9858 & tmp_ivl_9860;
  LPM_q_ivl_9864 <= tmp_ivl_9866 & tmp_ivl_9861;
  tmp_ivl_9869 <= z4(37);
  tmp_ivl_9870 <= new_AGEMA_signal_3141 & tmp_ivl_9869;
  LPM_q_ivl_9873 <= tmp_ivl_9875 & tmp_ivl_9870;
  new_AGEMA_signal_3328 <= tmp_ivl_9877(1);
  n3477 <= tmp_ivl_9877(0);
  tmp_ivl_9877 <= LPM_d0_ivl_9881(0 + 1 downto 0);
  tmp_ivl_9883 <= state_in_s1(285);
  tmp_ivl_9885 <= state_in_s0(285);
  tmp_ivl_9886 <= tmp_ivl_9883 & tmp_ivl_9885;
  LPM_q_ivl_9889 <= tmp_ivl_9891 & tmp_ivl_9886;
  tmp_ivl_9893 <= new_AGEMA_signal_3328 & n3477;
  LPM_q_ivl_9896 <= tmp_ivl_9898 & tmp_ivl_9893;
  new_AGEMA_signal_3618 <= tmp_ivl_9900(1);
  n3629 <= tmp_ivl_9900(0);
  tmp_ivl_9900 <= LPM_d0_ivl_9904(0 + 1 downto 0);
  tmp_ivl_9905 <= new_AGEMA_signal_3595 & n3836;
  LPM_q_ivl_9908 <= tmp_ivl_9910 & tmp_ivl_9905;
  tmp_ivl_9912 <= new_AGEMA_signal_3618 & n3629;
  LPM_q_ivl_9915 <= tmp_ivl_9917 & tmp_ivl_9912;
  new_AGEMA_signal_3905 <= tmp_ivl_9919(1);
  n3308 <= tmp_ivl_9919(0);
  tmp_ivl_9919 <= LPM_d0_ivl_9923(0 + 1 downto 0);
  tmp_ivl_9925 <= state_in_s1(246);
  tmp_ivl_9927 <= state_in_s0(246);
  tmp_ivl_9928 <= tmp_ivl_9925 & tmp_ivl_9927;
  LPM_q_ivl_9931 <= tmp_ivl_9933 & tmp_ivl_9928;
  tmp_ivl_9936 <= z4(14);
  tmp_ivl_9937 <= new_AGEMA_signal_3116 & tmp_ivl_9936;
  LPM_q_ivl_9940 <= tmp_ivl_9942 & tmp_ivl_9937;
  new_AGEMA_signal_3329 <= tmp_ivl_9944(1);
  n3598 <= tmp_ivl_9944(0);
  tmp_ivl_9944 <= LPM_d0_ivl_9948(0 + 1 downto 0);
  tmp_ivl_9950 <= state_in_s1(310);
  tmp_ivl_9952 <= state_in_s0(310);
  tmp_ivl_9953 <= tmp_ivl_9950 & tmp_ivl_9952;
  LPM_q_ivl_9956 <= tmp_ivl_9958 & tmp_ivl_9953;
  tmp_ivl_9960 <= new_AGEMA_signal_3329 & n3598;
  LPM_q_ivl_9963 <= tmp_ivl_9965 & tmp_ivl_9960;
  new_AGEMA_signal_3619 <= tmp_ivl_9967(1);
  n3377 <= tmp_ivl_9967(0);
  tmp_ivl_9967 <= LPM_d0_ivl_9971(0 + 1 downto 0);
  tmp_ivl_9972 <= new_AGEMA_signal_3905 & n3308;
  LPM_q_ivl_9975 <= tmp_ivl_9977 & tmp_ivl_9972;
  tmp_ivl_9979 <= new_AGEMA_signal_3619 & n3377;
  LPM_q_ivl_9982 <= tmp_ivl_9984 & tmp_ivl_9979;
  tmp_ivl_9986 <= tmp_ivl_9990(1);
  tmp_ivl_9988 <= tmp_ivl_9990(0);
  tmp_ivl_9990 <= LPM_d0_ivl_9994(0 + 1 downto 0);
  tmp_ivl_9996 <= state_in_s1(237);
  tmp_ivl_9998 <= state_in_s0(237);
  tmp_ivl_9999 <= tmp_ivl_9996 & tmp_ivl_9998;
  LPM_q_ivl_10002 <= '0' & tmp_ivl_9999;
  tmp_ivl_10007 <= z4(21);
  tmp_ivl_10008 <= new_AGEMA_signal_3124 & tmp_ivl_10007;
  LPM_q_ivl_10011 <= '0' & tmp_ivl_10008;
  new_AGEMA_signal_3330 <= tmp_ivl_10015(1);
  n3494 <= tmp_ivl_10015(0);
  tmp_ivl_10015 <= LPM_d0_ivl_10019(0 + 1 downto 0);
  tmp_ivl_10021 <= state_in_s1(301);
  tmp_ivl_10023 <= state_in_s0(301);
  tmp_ivl_10024 <= tmp_ivl_10021 & tmp_ivl_10023;
  LPM_q_ivl_10027 <= '0' & tmp_ivl_10024;
  tmp_ivl_10031 <= new_AGEMA_signal_3330 & n3494;
  LPM_q_ivl_10034 <= '0' & tmp_ivl_10031;
  new_AGEMA_signal_3620 <= tmp_ivl_10038(1);
  n3835 <= tmp_ivl_10038(0);
  tmp_ivl_10038 <= LPM_d0_ivl_10042(0 + 1 downto 0);
  tmp_ivl_10043 <= new_AGEMA_signal_3619 & n3377;
  LPM_q_ivl_10046 <= tmp_ivl_10048 & tmp_ivl_10043;
  tmp_ivl_10050 <= new_AGEMA_signal_3620 & n3835;
  LPM_q_ivl_10053 <= tmp_ivl_10055 & tmp_ivl_10050;
  new_AGEMA_signal_3906 <= tmp_ivl_10057(1);
  n3309 <= tmp_ivl_10057(0);
  tmp_ivl_10057 <= LPM_d0_ivl_10061(0 + 1 downto 0);
  tmp_ivl_10063 <= state_in_s1(207);
  tmp_ivl_10065 <= state_in_s0(207);
  tmp_ivl_10066 <= tmp_ivl_10063 & tmp_ivl_10065;
  LPM_q_ivl_10069 <= tmp_ivl_10071 & tmp_ivl_10066;
  tmp_ivl_10074 <= z4(55);
  tmp_ivl_10075 <= new_AGEMA_signal_3161 & tmp_ivl_10074;
  LPM_q_ivl_10078 <= tmp_ivl_10080 & tmp_ivl_10075;
  new_AGEMA_signal_3331 <= tmp_ivl_10082(1);
  n3394 <= tmp_ivl_10082(0);
  tmp_ivl_10082 <= LPM_d0_ivl_10086(0 + 1 downto 0);
  tmp_ivl_10088 <= state_in_s1(271);
  tmp_ivl_10090 <= state_in_s0(271);
  tmp_ivl_10091 <= tmp_ivl_10088 & tmp_ivl_10090;
  LPM_q_ivl_10094 <= tmp_ivl_10096 & tmp_ivl_10091;
  tmp_ivl_10098 <= new_AGEMA_signal_3331 & n3394;
  LPM_q_ivl_10101 <= tmp_ivl_10103 & tmp_ivl_10098;
  new_AGEMA_signal_3621 <= tmp_ivl_10105(1);
  n3510 <= tmp_ivl_10105(0);
  tmp_ivl_10105 <= LPM_d0_ivl_10109(0 + 1 downto 0);
  tmp_ivl_10110 <= new_AGEMA_signal_3906 & n3309;
  LPM_q_ivl_10113 <= tmp_ivl_10115 & tmp_ivl_10110;
  tmp_ivl_10117 <= new_AGEMA_signal_3621 & n3510;
  LPM_q_ivl_10120 <= tmp_ivl_10122 & tmp_ivl_10117;
  tmp_ivl_10124 <= tmp_ivl_10128(1);
  tmp_ivl_10126 <= tmp_ivl_10128(0);
  tmp_ivl_10128 <= LPM_d0_ivl_10132(0 + 1 downto 0);
  tmp_ivl_10134 <= z0(58);
  tmp_ivl_10135 <= new_AGEMA_signal_3249 & tmp_ivl_10134;
  LPM_q_ivl_10138 <= tmp_ivl_10140 & tmp_ivl_10135;
  tmp_ivl_10143 <= state_in_s1(2);
  tmp_ivl_10145 <= state_in_s0(2);
  tmp_ivl_10146 <= tmp_ivl_10143 & tmp_ivl_10145;
  LPM_q_ivl_10149 <= tmp_ivl_10151 & tmp_ivl_10146;
  new_AGEMA_signal_3332 <= tmp_ivl_10153(1);
  n3407 <= tmp_ivl_10153(0);
  tmp_ivl_10153 <= LPM_d0_ivl_10157(0 + 1 downto 0);
  tmp_ivl_10159 <= z1(58);
  tmp_ivl_10160 <= new_AGEMA_signal_3039 & tmp_ivl_10159;
  LPM_q_ivl_10163 <= tmp_ivl_10165 & tmp_ivl_10160;
  tmp_ivl_10167 <= new_AGEMA_signal_3332 & n3407;
  LPM_q_ivl_10170 <= tmp_ivl_10172 & tmp_ivl_10167;
  new_AGEMA_signal_3622 <= tmp_ivl_10174(1);
  n3311 <= tmp_ivl_10174(0);
  tmp_ivl_10174 <= LPM_d0_ivl_10178(0 + 1 downto 0);
  tmp_ivl_10179 <= new_AGEMA_signal_3622 & n3311;
  LPM_q_ivl_10182 <= tmp_ivl_10184 & tmp_ivl_10179;
  tmp_ivl_10186 <= new_AGEMA_signal_2657 & n3310;
  LPM_q_ivl_10189 <= tmp_ivl_10191 & tmp_ivl_10186;
  new_AGEMA_signal_3907 <= tmp_ivl_10193(1);
  n3542 <= tmp_ivl_10193(0);
  tmp_ivl_10193 <= LPM_d0_ivl_10197(0 + 1 downto 0);
  tmp_ivl_10199 <= z1(33);
  tmp_ivl_10200 <= new_AGEMA_signal_3014 & tmp_ivl_10199;
  LPM_q_ivl_10203 <= tmp_ivl_10205 & tmp_ivl_10200;
  tmp_ivl_10208 <= state_in_s1(281);
  tmp_ivl_10210 <= state_in_s0(281);
  tmp_ivl_10211 <= tmp_ivl_10208 & tmp_ivl_10210;
  LPM_q_ivl_10214 <= tmp_ivl_10216 & tmp_ivl_10211;
  new_AGEMA_signal_3333 <= tmp_ivl_10218(1);
  n3313 <= tmp_ivl_10218(0);
  tmp_ivl_10218 <= LPM_d0_ivl_10222(0 + 1 downto 0);
  tmp_ivl_10224 <= z0(33);
  tmp_ivl_10225 <= new_AGEMA_signal_3267 & tmp_ivl_10224;
  LPM_q_ivl_10228 <= tmp_ivl_10230 & tmp_ivl_10225;
  tmp_ivl_10233 <= state_in_s1(25);
  tmp_ivl_10235 <= state_in_s0(25);
  tmp_ivl_10236 <= tmp_ivl_10233 & tmp_ivl_10235;
  LPM_q_ivl_10239 <= tmp_ivl_10241 & tmp_ivl_10236;
  new_AGEMA_signal_3334 <= tmp_ivl_10243(1);
  n3614 <= tmp_ivl_10243(0);
  tmp_ivl_10243 <= LPM_d0_ivl_10247(0 + 1 downto 0);
  tmp_ivl_10249 <= state_in_s1(89);
  tmp_ivl_10251 <= state_in_s0(89);
  tmp_ivl_10252 <= tmp_ivl_10249 & tmp_ivl_10251;
  LPM_q_ivl_10255 <= tmp_ivl_10257 & tmp_ivl_10252;
  tmp_ivl_10259 <= new_AGEMA_signal_3334 & n3614;
  LPM_q_ivl_10262 <= tmp_ivl_10264 & tmp_ivl_10259;
  new_AGEMA_signal_3623 <= tmp_ivl_10266(1);
  n3312 <= tmp_ivl_10266(0);
  tmp_ivl_10266 <= LPM_d0_ivl_10270(0 + 1 downto 0);
  tmp_ivl_10271 <= new_AGEMA_signal_3333 & n3313;
  LPM_q_ivl_10274 <= tmp_ivl_10276 & tmp_ivl_10271;
  tmp_ivl_10278 <= new_AGEMA_signal_3623 & n3312;
  LPM_q_ivl_10281 <= tmp_ivl_10283 & tmp_ivl_10278;
  new_AGEMA_signal_3908 <= tmp_ivl_10285(1);
  n3447 <= tmp_ivl_10285(0);
  tmp_ivl_10285 <= LPM_d0_ivl_10289(0 + 1 downto 0);
  tmp_ivl_10290 <= new_AGEMA_signal_3907 & n3542;
  LPM_q_ivl_10293 <= tmp_ivl_10295 & tmp_ivl_10290;
  tmp_ivl_10297 <= new_AGEMA_signal_3908 & n3447;
  LPM_q_ivl_10300 <= tmp_ivl_10302 & tmp_ivl_10297;
  new_AGEMA_signal_4220 <= tmp_ivl_10304(1);
  n3316 <= tmp_ivl_10304(0);
  tmp_ivl_10304 <= LPM_d0_ivl_10308(0 + 1 downto 0);
  tmp_ivl_10310 <= z1(55);
  tmp_ivl_10311 <= new_AGEMA_signal_3036 & tmp_ivl_10310;
  LPM_q_ivl_10314 <= tmp_ivl_10316 & tmp_ivl_10311;
  tmp_ivl_10319 <= state_in_s1(271);
  tmp_ivl_10321 <= state_in_s0(271);
  tmp_ivl_10322 <= tmp_ivl_10319 & tmp_ivl_10321;
  LPM_q_ivl_10325 <= tmp_ivl_10327 & tmp_ivl_10322;
  new_AGEMA_signal_3335 <= tmp_ivl_10329(1);
  n3315 <= tmp_ivl_10329(0);
  tmp_ivl_10329 <= LPM_d0_ivl_10333(0 + 1 downto 0);
  tmp_ivl_10335 <= z0(55);
  tmp_ivl_10336 <= new_AGEMA_signal_3253 & tmp_ivl_10335;
  LPM_q_ivl_10339 <= tmp_ivl_10341 & tmp_ivl_10336;
  tmp_ivl_10344 <= state_in_s1(15);
  tmp_ivl_10346 <= state_in_s0(15);
  tmp_ivl_10347 <= tmp_ivl_10344 & tmp_ivl_10346;
  LPM_q_ivl_10350 <= tmp_ivl_10352 & tmp_ivl_10347;
  new_AGEMA_signal_3336 <= tmp_ivl_10354(1);
  n3395 <= tmp_ivl_10354(0);
  tmp_ivl_10354 <= LPM_d0_ivl_10358(0 + 1 downto 0);
  tmp_ivl_10360 <= state_in_s1(79);
  tmp_ivl_10362 <= state_in_s0(79);
  tmp_ivl_10363 <= tmp_ivl_10360 & tmp_ivl_10362;
  LPM_q_ivl_10366 <= tmp_ivl_10368 & tmp_ivl_10363;
  tmp_ivl_10370 <= new_AGEMA_signal_3336 & n3395;
  LPM_q_ivl_10373 <= tmp_ivl_10375 & tmp_ivl_10370;
  new_AGEMA_signal_3624 <= tmp_ivl_10377(1);
  n3314 <= tmp_ivl_10377(0);
  tmp_ivl_10377 <= LPM_d0_ivl_10381(0 + 1 downto 0);
  tmp_ivl_10382 <= new_AGEMA_signal_3335 & n3315;
  LPM_q_ivl_10385 <= tmp_ivl_10387 & tmp_ivl_10382;
  tmp_ivl_10389 <= new_AGEMA_signal_3624 & n3314;
  LPM_q_ivl_10392 <= tmp_ivl_10394 & tmp_ivl_10389;
  new_AGEMA_signal_3909 <= tmp_ivl_10396(1);
  n3433 <= tmp_ivl_10396(0);
  tmp_ivl_10396 <= LPM_d0_ivl_10400(0 + 1 downto 0);
  tmp_ivl_10401 <= new_AGEMA_signal_4220 & n3316;
  LPM_q_ivl_10404 <= tmp_ivl_10406 & tmp_ivl_10401;
  tmp_ivl_10408 <= new_AGEMA_signal_3909 & n3433;
  LPM_q_ivl_10411 <= tmp_ivl_10413 & tmp_ivl_10408;
  tmp_ivl_10415 <= tmp_ivl_10419(1);
  tmp_ivl_10417 <= tmp_ivl_10419(0);
  tmp_ivl_10419 <= LPM_d0_ivl_10423(0 + 1 downto 0);
  tmp_ivl_10425 <= z0(59);
  tmp_ivl_10426 <= new_AGEMA_signal_3247 & tmp_ivl_10425;
  LPM_q_ivl_10429 <= tmp_ivl_10431 & tmp_ivl_10426;
  tmp_ivl_10434 <= state_in_s1(3);
  tmp_ivl_10436 <= state_in_s0(3);
  tmp_ivl_10437 <= tmp_ivl_10434 & tmp_ivl_10436;
  LPM_q_ivl_10440 <= tmp_ivl_10442 & tmp_ivl_10437;
  new_AGEMA_signal_3337 <= tmp_ivl_10444(1);
  n3597 <= tmp_ivl_10444(0);
  tmp_ivl_10444 <= LPM_d0_ivl_10448(0 + 1 downto 0);
  tmp_ivl_10450 <= z1(59);
  tmp_ivl_10451 <= new_AGEMA_signal_3040 & tmp_ivl_10450;
  LPM_q_ivl_10454 <= tmp_ivl_10456 & tmp_ivl_10451;
  tmp_ivl_10458 <= new_AGEMA_signal_3337 & n3597;
  LPM_q_ivl_10461 <= tmp_ivl_10463 & tmp_ivl_10458;
  new_AGEMA_signal_3625 <= tmp_ivl_10465(1);
  n3318 <= tmp_ivl_10465(0);
  tmp_ivl_10465 <= LPM_d0_ivl_10469(0 + 1 downto 0);
  tmp_ivl_10470 <= new_AGEMA_signal_3625 & n3318;
  LPM_q_ivl_10473 <= tmp_ivl_10475 & tmp_ivl_10470;
  tmp_ivl_10477 <= new_AGEMA_signal_2659 & n3317;
  LPM_q_ivl_10480 <= tmp_ivl_10482 & tmp_ivl_10477;
  new_AGEMA_signal_3910 <= tmp_ivl_10484(1);
  n3572 <= tmp_ivl_10484(0);
  tmp_ivl_10484 <= LPM_d0_ivl_10488(0 + 1 downto 0);
  tmp_ivl_10490 <= z1(34);
  tmp_ivl_10491 <= new_AGEMA_signal_3015 & tmp_ivl_10490;
  LPM_q_ivl_10494 <= tmp_ivl_10496 & tmp_ivl_10491;
  tmp_ivl_10499 <= state_in_s1(282);
  tmp_ivl_10501 <= state_in_s0(282);
  tmp_ivl_10502 <= tmp_ivl_10499 & tmp_ivl_10501;
  LPM_q_ivl_10505 <= tmp_ivl_10507 & tmp_ivl_10502;
  new_AGEMA_signal_3338 <= tmp_ivl_10509(1);
  n3320 <= tmp_ivl_10509(0);
  tmp_ivl_10509 <= LPM_d0_ivl_10513(0 + 1 downto 0);
  tmp_ivl_10515 <= z0(34);
  tmp_ivl_10516 <= new_AGEMA_signal_3265 & tmp_ivl_10515;
  LPM_q_ivl_10519 <= tmp_ivl_10521 & tmp_ivl_10516;
  tmp_ivl_10524 <= state_in_s1(26);
  tmp_ivl_10526 <= state_in_s0(26);
  tmp_ivl_10527 <= tmp_ivl_10524 & tmp_ivl_10526;
  LPM_q_ivl_10530 <= tmp_ivl_10532 & tmp_ivl_10527;
  new_AGEMA_signal_3339 <= tmp_ivl_10534(1);
  n3569 <= tmp_ivl_10534(0);
  tmp_ivl_10534 <= LPM_d0_ivl_10538(0 + 1 downto 0);
  tmp_ivl_10540 <= state_in_s1(90);
  tmp_ivl_10542 <= state_in_s0(90);
  tmp_ivl_10543 <= tmp_ivl_10540 & tmp_ivl_10542;
  LPM_q_ivl_10546 <= tmp_ivl_10548 & tmp_ivl_10543;
  tmp_ivl_10550 <= new_AGEMA_signal_3339 & n3569;
  LPM_q_ivl_10553 <= tmp_ivl_10555 & tmp_ivl_10550;
  new_AGEMA_signal_3626 <= tmp_ivl_10557(1);
  n3319 <= tmp_ivl_10557(0);
  tmp_ivl_10557 <= LPM_d0_ivl_10561(0 + 1 downto 0);
  tmp_ivl_10562 <= new_AGEMA_signal_3338 & n3320;
  LPM_q_ivl_10565 <= tmp_ivl_10567 & tmp_ivl_10562;
  tmp_ivl_10569 <= new_AGEMA_signal_3626 & n3319;
  LPM_q_ivl_10572 <= tmp_ivl_10574 & tmp_ivl_10569;
  new_AGEMA_signal_3911 <= tmp_ivl_10576(1);
  n3502 <= tmp_ivl_10576(0);
  tmp_ivl_10576 <= LPM_d0_ivl_10580(0 + 1 downto 0);
  tmp_ivl_10581 <= new_AGEMA_signal_3910 & n3572;
  LPM_q_ivl_10584 <= tmp_ivl_10586 & tmp_ivl_10581;
  tmp_ivl_10588 <= new_AGEMA_signal_3911 & n3502;
  LPM_q_ivl_10591 <= tmp_ivl_10593 & tmp_ivl_10588;
  new_AGEMA_signal_4221 <= tmp_ivl_10595(1);
  n3323 <= tmp_ivl_10595(0);
  tmp_ivl_10595 <= LPM_d0_ivl_10599(0 + 1 downto 0);
  tmp_ivl_10601 <= z1(56);
  tmp_ivl_10602 <= new_AGEMA_signal_3037 & tmp_ivl_10601;
  LPM_q_ivl_10605 <= tmp_ivl_10607 & tmp_ivl_10602;
  tmp_ivl_10610 <= state_in_s1(256);
  tmp_ivl_10612 <= state_in_s0(256);
  tmp_ivl_10613 <= tmp_ivl_10610 & tmp_ivl_10612;
  LPM_q_ivl_10616 <= tmp_ivl_10618 & tmp_ivl_10613;
  new_AGEMA_signal_3340 <= tmp_ivl_10620(1);
  n3322 <= tmp_ivl_10620(0);
  tmp_ivl_10620 <= LPM_d0_ivl_10624(0 + 1 downto 0);
  tmp_ivl_10626 <= z0(56);
  tmp_ivl_10627 <= new_AGEMA_signal_3252 & tmp_ivl_10626;
  LPM_q_ivl_10630 <= tmp_ivl_10632 & tmp_ivl_10627;
  tmp_ivl_10635 <= state_in_s1(0);
  tmp_ivl_10637 <= state_in_s0(0);
  tmp_ivl_10638 <= tmp_ivl_10635 & tmp_ivl_10637;
  LPM_q_ivl_10641 <= tmp_ivl_10643 & tmp_ivl_10638;
  new_AGEMA_signal_3341 <= tmp_ivl_10645(1);
  n3442 <= tmp_ivl_10645(0);
  tmp_ivl_10645 <= LPM_d0_ivl_10649(0 + 1 downto 0);
  tmp_ivl_10651 <= state_in_s1(64);
  tmp_ivl_10653 <= state_in_s0(64);
  tmp_ivl_10654 <= tmp_ivl_10651 & tmp_ivl_10653;
  LPM_q_ivl_10657 <= tmp_ivl_10659 & tmp_ivl_10654;
  tmp_ivl_10661 <= new_AGEMA_signal_3341 & n3442;
  LPM_q_ivl_10664 <= tmp_ivl_10666 & tmp_ivl_10661;
  new_AGEMA_signal_3627 <= tmp_ivl_10668(1);
  n3321 <= tmp_ivl_10668(0);
  tmp_ivl_10668 <= LPM_d0_ivl_10672(0 + 1 downto 0);
  tmp_ivl_10673 <= new_AGEMA_signal_3340 & n3322;
  LPM_q_ivl_10676 <= tmp_ivl_10678 & tmp_ivl_10673;
  tmp_ivl_10680 <= new_AGEMA_signal_3627 & n3321;
  LPM_q_ivl_10683 <= tmp_ivl_10685 & tmp_ivl_10680;
  new_AGEMA_signal_3912 <= tmp_ivl_10687(1);
  n3464 <= tmp_ivl_10687(0);
  tmp_ivl_10687 <= LPM_d0_ivl_10691(0 + 1 downto 0);
  tmp_ivl_10692 <= new_AGEMA_signal_4221 & n3323;
  LPM_q_ivl_10695 <= tmp_ivl_10697 & tmp_ivl_10692;
  tmp_ivl_10699 <= new_AGEMA_signal_3912 & n3464;
  LPM_q_ivl_10702 <= tmp_ivl_10704 & tmp_ivl_10699;
  tmp_ivl_10706 <= tmp_ivl_10710(1);
  tmp_ivl_10708 <= tmp_ivl_10710(0);
  tmp_ivl_10710 <= LPM_d0_ivl_10714(0 + 1 downto 0);
  tmp_ivl_10715 <= new_AGEMA_signal_3586 & n3664;
  LPM_q_ivl_10718 <= tmp_ivl_10720 & tmp_ivl_10715;
  tmp_ivl_10722 <= new_AGEMA_signal_3598 & n3925;
  LPM_q_ivl_10725 <= tmp_ivl_10727 & tmp_ivl_10722;
  new_AGEMA_signal_3913 <= tmp_ivl_10729(1);
  n3324 <= tmp_ivl_10729(0);
  tmp_ivl_10729 <= LPM_d0_ivl_10733(0 + 1 downto 0);
  tmp_ivl_10735 <= state_in_s1(222);
  tmp_ivl_10737 <= state_in_s0(222);
  tmp_ivl_10738 <= tmp_ivl_10735 & tmp_ivl_10737;
  LPM_q_ivl_10741 <= tmp_ivl_10743 & tmp_ivl_10738;
  tmp_ivl_10746 <= z4(38);
  tmp_ivl_10747 <= new_AGEMA_signal_3142 & tmp_ivl_10746;
  LPM_q_ivl_10750 <= tmp_ivl_10752 & tmp_ivl_10747;
  new_AGEMA_signal_3342 <= tmp_ivl_10754(1);
  n3353 <= tmp_ivl_10754(0);
  tmp_ivl_10754 <= LPM_d0_ivl_10758(0 + 1 downto 0);
  tmp_ivl_10760 <= state_in_s1(286);
  tmp_ivl_10762 <= state_in_s0(286);
  tmp_ivl_10763 <= tmp_ivl_10760 & tmp_ivl_10762;
  LPM_q_ivl_10766 <= tmp_ivl_10768 & tmp_ivl_10763;
  tmp_ivl_10770 <= new_AGEMA_signal_3342 & n3353;
  LPM_q_ivl_10773 <= tmp_ivl_10775 & tmp_ivl_10770;
  new_AGEMA_signal_3628 <= tmp_ivl_10777(1);
  n3453 <= tmp_ivl_10777(0);
  tmp_ivl_10777 <= LPM_d0_ivl_10781(0 + 1 downto 0);
  tmp_ivl_10782 <= new_AGEMA_signal_3913 & n3324;
  LPM_q_ivl_10785 <= tmp_ivl_10787 & tmp_ivl_10782;
  tmp_ivl_10789 <= new_AGEMA_signal_3628 & n3453;
  LPM_q_ivl_10792 <= tmp_ivl_10794 & tmp_ivl_10789;
  tmp_ivl_10796 <= tmp_ivl_10800(1);
  tmp_ivl_10798 <= tmp_ivl_10800(0);
  tmp_ivl_10800 <= LPM_d0_ivl_10804(0 + 1 downto 0);
  tmp_ivl_10805 <= new_AGEMA_signal_3588 & n3663;
  LPM_q_ivl_10808 <= tmp_ivl_10810 & tmp_ivl_10805;
  tmp_ivl_10812 <= new_AGEMA_signal_3628 & n3453;
  LPM_q_ivl_10815 <= tmp_ivl_10817 & tmp_ivl_10812;
  new_AGEMA_signal_3914 <= tmp_ivl_10819(1);
  n3325 <= tmp_ivl_10819(0);
  tmp_ivl_10819 <= LPM_d0_ivl_10823(0 + 1 downto 0);
  tmp_ivl_10825 <= state_in_s1(231);
  tmp_ivl_10827 <= state_in_s0(231);
  tmp_ivl_10828 <= tmp_ivl_10825 & tmp_ivl_10827;
  LPM_q_ivl_10831 <= tmp_ivl_10833 & tmp_ivl_10828;
  tmp_ivl_10836 <= z4(31);
  tmp_ivl_10837 <= new_AGEMA_signal_3135 & tmp_ivl_10836;
  LPM_q_ivl_10840 <= tmp_ivl_10842 & tmp_ivl_10837;
  new_AGEMA_signal_3343 <= tmp_ivl_10844(1);
  n3551 <= tmp_ivl_10844(0);
  tmp_ivl_10844 <= LPM_d0_ivl_10848(0 + 1 downto 0);
  tmp_ivl_10850 <= state_in_s1(295);
  tmp_ivl_10852 <= state_in_s0(295);
  tmp_ivl_10853 <= tmp_ivl_10850 & tmp_ivl_10852;
  LPM_q_ivl_10856 <= tmp_ivl_10858 & tmp_ivl_10853;
  tmp_ivl_10860 <= new_AGEMA_signal_3343 & n3551;
  LPM_q_ivl_10863 <= tmp_ivl_10865 & tmp_ivl_10860;
  new_AGEMA_signal_3629 <= tmp_ivl_10867(1);
  n3456 <= tmp_ivl_10867(0);
  tmp_ivl_10867 <= LPM_d0_ivl_10871(0 + 1 downto 0);
  tmp_ivl_10872 <= new_AGEMA_signal_3914 & n3325;
  LPM_q_ivl_10875 <= tmp_ivl_10877 & tmp_ivl_10872;
  tmp_ivl_10879 <= new_AGEMA_signal_3629 & n3456;
  LPM_q_ivl_10882 <= tmp_ivl_10884 & tmp_ivl_10879;
  tmp_ivl_10886 <= tmp_ivl_10890(1);
  tmp_ivl_10888 <= tmp_ivl_10890(0);
  tmp_ivl_10890 <= LPM_d0_ivl_10894(0 + 1 downto 0);
  tmp_ivl_10896 <= state_in_s1(193);
  tmp_ivl_10898 <= state_in_s0(193);
  tmp_ivl_10899 <= tmp_ivl_10896 & tmp_ivl_10898;
  LPM_q_ivl_10902 <= tmp_ivl_10904 & tmp_ivl_10899;
  tmp_ivl_10907 <= z4(57);
  tmp_ivl_10908 <= new_AGEMA_signal_3163 & tmp_ivl_10907;
  LPM_q_ivl_10911 <= tmp_ivl_10913 & tmp_ivl_10908;
  new_AGEMA_signal_3344 <= tmp_ivl_10915(1);
  n3496 <= tmp_ivl_10915(0);
  tmp_ivl_10915 <= LPM_d0_ivl_10919(0 + 1 downto 0);
  tmp_ivl_10921 <= state_in_s1(257);
  tmp_ivl_10923 <= state_in_s0(257);
  tmp_ivl_10924 <= tmp_ivl_10921 & tmp_ivl_10923;
  LPM_q_ivl_10927 <= tmp_ivl_10929 & tmp_ivl_10924;
  tmp_ivl_10931 <= new_AGEMA_signal_3344 & n3496;
  LPM_q_ivl_10934 <= tmp_ivl_10936 & tmp_ivl_10931;
  new_AGEMA_signal_3630 <= tmp_ivl_10938(1);
  n3726 <= tmp_ivl_10938(0);
  tmp_ivl_10938 <= LPM_d0_ivl_10942(0 + 1 downto 0);
  tmp_ivl_10943 <= new_AGEMA_signal_3615 & n3422;
  LPM_q_ivl_10946 <= tmp_ivl_10948 & tmp_ivl_10943;
  tmp_ivl_10950 <= new_AGEMA_signal_3630 & n3726;
  LPM_q_ivl_10953 <= tmp_ivl_10955 & tmp_ivl_10950;
  new_AGEMA_signal_3915 <= tmp_ivl_10957(1);
  n3326 <= tmp_ivl_10957(0);
  tmp_ivl_10957 <= LPM_d0_ivl_10961(0 + 1 downto 0);
  tmp_ivl_10963 <= state_in_s1(248);
  tmp_ivl_10965 <= state_in_s0(248);
  tmp_ivl_10966 <= tmp_ivl_10963 & tmp_ivl_10965;
  LPM_q_ivl_10969 <= tmp_ivl_10971 & tmp_ivl_10966;
  tmp_ivl_10974 <= z4(0);
  tmp_ivl_10975 <= new_AGEMA_signal_3111 & tmp_ivl_10974;
  LPM_q_ivl_10978 <= tmp_ivl_10980 & tmp_ivl_10975;
  new_AGEMA_signal_3345 <= tmp_ivl_10982(1);
  n3634 <= tmp_ivl_10982(0);
  tmp_ivl_10982 <= LPM_d0_ivl_10986(0 + 1 downto 0);
  tmp_ivl_10988 <= state_in_s1(312);
  tmp_ivl_10990 <= state_in_s0(312);
  tmp_ivl_10991 <= tmp_ivl_10988 & tmp_ivl_10990;
  LPM_q_ivl_10994 <= tmp_ivl_10996 & tmp_ivl_10991;
  tmp_ivl_10998 <= new_AGEMA_signal_3345 & n3634;
  LPM_q_ivl_11001 <= tmp_ivl_11003 & tmp_ivl_10998;
  new_AGEMA_signal_3631 <= tmp_ivl_11005(1);
  n3631 <= tmp_ivl_11005(0);
  tmp_ivl_11005 <= LPM_d0_ivl_11009(0 + 1 downto 0);
  tmp_ivl_11010 <= new_AGEMA_signal_3915 & n3326;
  LPM_q_ivl_11013 <= tmp_ivl_11015 & tmp_ivl_11010;
  tmp_ivl_11017 <= new_AGEMA_signal_3631 & n3631;
  LPM_q_ivl_11020 <= tmp_ivl_11022 & tmp_ivl_11017;
  tmp_ivl_11024 <= tmp_ivl_11028(1);
  tmp_ivl_11026 <= tmp_ivl_11028(0);
  tmp_ivl_11028 <= LPM_d0_ivl_11032(0 + 1 downto 0);
  tmp_ivl_11034 <= z1(60);
  tmp_ivl_11035 <= new_AGEMA_signal_3041 & tmp_ivl_11034;
  LPM_q_ivl_11038 <= tmp_ivl_11040 & tmp_ivl_11035;
  tmp_ivl_11043 <= state_in_s1(260);
  tmp_ivl_11045 <= state_in_s0(260);
  tmp_ivl_11046 <= tmp_ivl_11043 & tmp_ivl_11045;
  LPM_q_ivl_11049 <= tmp_ivl_11051 & tmp_ivl_11046;
  new_AGEMA_signal_3346 <= tmp_ivl_11053(1);
  n3328 <= tmp_ivl_11053(0);
  tmp_ivl_11053 <= LPM_d0_ivl_11057(0 + 1 downto 0);
  tmp_ivl_11059 <= z0(60);
  tmp_ivl_11060 <= new_AGEMA_signal_3244 & tmp_ivl_11059;
  LPM_q_ivl_11063 <= tmp_ivl_11065 & tmp_ivl_11060;
  tmp_ivl_11068 <= state_in_s1(4);
  tmp_ivl_11070 <= state_in_s0(4);
  tmp_ivl_11071 <= tmp_ivl_11068 & tmp_ivl_11070;
  LPM_q_ivl_11074 <= tmp_ivl_11076 & tmp_ivl_11071;
  new_AGEMA_signal_3347 <= tmp_ivl_11078(1);
  n3486 <= tmp_ivl_11078(0);
  tmp_ivl_11078 <= LPM_d0_ivl_11082(0 + 1 downto 0);
  tmp_ivl_11084 <= state_in_s1(68);
  tmp_ivl_11086 <= state_in_s0(68);
  tmp_ivl_11087 <= tmp_ivl_11084 & tmp_ivl_11086;
  LPM_q_ivl_11090 <= tmp_ivl_11092 & tmp_ivl_11087;
  tmp_ivl_11094 <= new_AGEMA_signal_3347 & n3486;
  LPM_q_ivl_11097 <= tmp_ivl_11099 & tmp_ivl_11094;
  new_AGEMA_signal_3632 <= tmp_ivl_11101(1);
  n3327 <= tmp_ivl_11101(0);
  tmp_ivl_11101 <= LPM_d0_ivl_11105(0 + 1 downto 0);
  tmp_ivl_11106 <= new_AGEMA_signal_3346 & n3328;
  LPM_q_ivl_11109 <= tmp_ivl_11111 & tmp_ivl_11106;
  tmp_ivl_11113 <= new_AGEMA_signal_3632 & n3327;
  LPM_q_ivl_11116 <= tmp_ivl_11118 & tmp_ivl_11113;
  new_AGEMA_signal_3916 <= tmp_ivl_11120(1);
  n3586 <= tmp_ivl_11120(0);
  tmp_ivl_11120 <= LPM_d0_ivl_11124(0 + 1 downto 0);
  tmp_ivl_11126 <= z0(57);
  tmp_ivl_11127 <= new_AGEMA_signal_3251 & tmp_ivl_11126;
  LPM_q_ivl_11130 <= tmp_ivl_11132 & tmp_ivl_11127;
  tmp_ivl_11135 <= state_in_s1(1);
  tmp_ivl_11137 <= state_in_s0(1);
  tmp_ivl_11138 <= tmp_ivl_11135 & tmp_ivl_11137;
  LPM_q_ivl_11141 <= tmp_ivl_11143 & tmp_ivl_11138;
  new_AGEMA_signal_3348 <= tmp_ivl_11145(1);
  n3497 <= tmp_ivl_11145(0);
  tmp_ivl_11145 <= LPM_d0_ivl_11149(0 + 1 downto 0);
  tmp_ivl_11151 <= z1(57);
  tmp_ivl_11152 <= new_AGEMA_signal_3038 & tmp_ivl_11151;
  LPM_q_ivl_11155 <= tmp_ivl_11157 & tmp_ivl_11152;
  tmp_ivl_11159 <= new_AGEMA_signal_3348 & n3497;
  LPM_q_ivl_11162 <= tmp_ivl_11164 & tmp_ivl_11159;
  new_AGEMA_signal_3633 <= tmp_ivl_11166(1);
  n3330 <= tmp_ivl_11166(0);
  tmp_ivl_11166 <= LPM_d0_ivl_11170(0 + 1 downto 0);
  tmp_ivl_11171 <= new_AGEMA_signal_3633 & n3330;
  LPM_q_ivl_11174 <= tmp_ivl_11176 & tmp_ivl_11171;
  tmp_ivl_11178 <= new_AGEMA_signal_2661 & n3329;
  LPM_q_ivl_11181 <= tmp_ivl_11183 & tmp_ivl_11178;
  new_AGEMA_signal_3917 <= tmp_ivl_11185(1);
  n3515 <= tmp_ivl_11185(0);
  tmp_ivl_11185 <= LPM_d0_ivl_11189(0 + 1 downto 0);
  tmp_ivl_11190 <= new_AGEMA_signal_3916 & n3586;
  LPM_q_ivl_11193 <= tmp_ivl_11195 & tmp_ivl_11190;
  tmp_ivl_11197 <= new_AGEMA_signal_3917 & n3515;
  LPM_q_ivl_11200 <= tmp_ivl_11202 & tmp_ivl_11197;
  new_AGEMA_signal_4225 <= tmp_ivl_11204(1);
  n3333 <= tmp_ivl_11204(0);
  tmp_ivl_11204 <= LPM_d0_ivl_11208(0 + 1 downto 0);
  tmp_ivl_11210 <= z1(35);
  tmp_ivl_11211 <= new_AGEMA_signal_3016 & tmp_ivl_11210;
  LPM_q_ivl_11214 <= tmp_ivl_11216 & tmp_ivl_11211;
  tmp_ivl_11219 <= state_in_s1(283);
  tmp_ivl_11221 <= state_in_s0(283);
  tmp_ivl_11222 <= tmp_ivl_11219 & tmp_ivl_11221;
  LPM_q_ivl_11225 <= tmp_ivl_11227 & tmp_ivl_11222;
  new_AGEMA_signal_3349 <= tmp_ivl_11229(1);
  n3332 <= tmp_ivl_11229(0);
  tmp_ivl_11229 <= LPM_d0_ivl_11233(0 + 1 downto 0);
  tmp_ivl_11235 <= z0(35);
  tmp_ivl_11236 <= new_AGEMA_signal_3263 & tmp_ivl_11235;
  LPM_q_ivl_11239 <= tmp_ivl_11241 & tmp_ivl_11236;
  tmp_ivl_11244 <= state_in_s1(27);
  tmp_ivl_11246 <= state_in_s0(27);
  tmp_ivl_11247 <= tmp_ivl_11244 & tmp_ivl_11246;
  LPM_q_ivl_11250 <= tmp_ivl_11252 & tmp_ivl_11247;
  new_AGEMA_signal_3350 <= tmp_ivl_11254(1);
  n3581 <= tmp_ivl_11254(0);
  tmp_ivl_11254 <= LPM_d0_ivl_11258(0 + 1 downto 0);
  tmp_ivl_11260 <= state_in_s1(91);
  tmp_ivl_11262 <= state_in_s0(91);
  tmp_ivl_11263 <= tmp_ivl_11260 & tmp_ivl_11262;
  LPM_q_ivl_11266 <= tmp_ivl_11268 & tmp_ivl_11263;
  tmp_ivl_11270 <= new_AGEMA_signal_3350 & n3581;
  LPM_q_ivl_11273 <= tmp_ivl_11275 & tmp_ivl_11270;
  new_AGEMA_signal_3634 <= tmp_ivl_11277(1);
  n3331 <= tmp_ivl_11277(0);
  tmp_ivl_11277 <= LPM_d0_ivl_11281(0 + 1 downto 0);
  tmp_ivl_11282 <= new_AGEMA_signal_3349 & n3332;
  LPM_q_ivl_11285 <= tmp_ivl_11287 & tmp_ivl_11282;
  tmp_ivl_11289 <= new_AGEMA_signal_3634 & n3331;
  LPM_q_ivl_11292 <= tmp_ivl_11294 & tmp_ivl_11289;
  new_AGEMA_signal_3918 <= tmp_ivl_11296(1);
  n3412 <= tmp_ivl_11296(0);
  tmp_ivl_11296 <= LPM_d0_ivl_11300(0 + 1 downto 0);
  tmp_ivl_11301 <= new_AGEMA_signal_4225 & n3333;
  LPM_q_ivl_11304 <= tmp_ivl_11306 & tmp_ivl_11301;
  tmp_ivl_11308 <= new_AGEMA_signal_3918 & n3412;
  LPM_q_ivl_11311 <= tmp_ivl_11313 & tmp_ivl_11308;
  tmp_ivl_11315 <= tmp_ivl_11319(1);
  tmp_ivl_11317 <= tmp_ivl_11319(0);
  tmp_ivl_11319 <= LPM_d0_ivl_11323(0 + 1 downto 0);
  tmp_ivl_11325 <= z1(21);
  tmp_ivl_11326 <= new_AGEMA_signal_3002 & tmp_ivl_11325;
  LPM_q_ivl_11329 <= tmp_ivl_11331 & tmp_ivl_11326;
  tmp_ivl_11334 <= state_in_s1(301);
  tmp_ivl_11336 <= state_in_s0(301);
  tmp_ivl_11337 <= tmp_ivl_11334 & tmp_ivl_11336;
  LPM_q_ivl_11340 <= tmp_ivl_11342 & tmp_ivl_11337;
  new_AGEMA_signal_3351 <= tmp_ivl_11344(1);
  n3335 <= tmp_ivl_11344(0);
  tmp_ivl_11344 <= LPM_d0_ivl_11348(0 + 1 downto 0);
  tmp_ivl_11350 <= z0(21);
  tmp_ivl_11351 <= new_AGEMA_signal_3245 & tmp_ivl_11350;
  LPM_q_ivl_11354 <= tmp_ivl_11356 & tmp_ivl_11351;
  tmp_ivl_11359 <= state_in_s1(45);
  tmp_ivl_11361 <= state_in_s0(45);
  tmp_ivl_11362 <= tmp_ivl_11359 & tmp_ivl_11361;
  LPM_q_ivl_11365 <= tmp_ivl_11367 & tmp_ivl_11362;
  new_AGEMA_signal_3352 <= tmp_ivl_11369(1);
  n3495 <= tmp_ivl_11369(0);
  tmp_ivl_11369 <= LPM_d0_ivl_11373(0 + 1 downto 0);
  tmp_ivl_11375 <= state_in_s1(109);
  tmp_ivl_11377 <= state_in_s0(109);
  tmp_ivl_11378 <= tmp_ivl_11375 & tmp_ivl_11377;
  LPM_q_ivl_11381 <= tmp_ivl_11383 & tmp_ivl_11378;
  tmp_ivl_11385 <= new_AGEMA_signal_3352 & n3495;
  LPM_q_ivl_11388 <= tmp_ivl_11390 & tmp_ivl_11385;
  new_AGEMA_signal_3635 <= tmp_ivl_11392(1);
  n3334 <= tmp_ivl_11392(0);
  tmp_ivl_11392 <= LPM_d0_ivl_11396(0 + 1 downto 0);
  tmp_ivl_11397 <= new_AGEMA_signal_3351 & n3335;
  LPM_q_ivl_11400 <= tmp_ivl_11402 & tmp_ivl_11397;
  tmp_ivl_11404 <= new_AGEMA_signal_3635 & n3334;
  LPM_q_ivl_11407 <= tmp_ivl_11409 & tmp_ivl_11404;
  new_AGEMA_signal_3919 <= tmp_ivl_11411(1);
  n3853 <= tmp_ivl_11411(0);
  tmp_ivl_11411 <= LPM_d0_ivl_11415(0 + 1 downto 0);
  tmp_ivl_11416 <= new_AGEMA_signal_3916 & n3586;
  LPM_q_ivl_11419 <= tmp_ivl_11421 & tmp_ivl_11416;
  tmp_ivl_11423 <= new_AGEMA_signal_3919 & n3853;
  LPM_q_ivl_11426 <= tmp_ivl_11428 & tmp_ivl_11423;
  new_AGEMA_signal_4226 <= tmp_ivl_11430(1);
  n3338 <= tmp_ivl_11430(0);
  tmp_ivl_11430 <= LPM_d0_ivl_11434(0 + 1 downto 0);
  tmp_ivl_11436 <= z0(18);
  tmp_ivl_11437 <= new_AGEMA_signal_3246 & tmp_ivl_11436;
  LPM_q_ivl_11440 <= tmp_ivl_11442 & tmp_ivl_11437;
  tmp_ivl_11445 <= state_in_s1(42);
  tmp_ivl_11447 <= state_in_s0(42);
  tmp_ivl_11448 <= tmp_ivl_11445 & tmp_ivl_11447;
  LPM_q_ivl_11451 <= tmp_ivl_11453 & tmp_ivl_11448;
  new_AGEMA_signal_3353 <= tmp_ivl_11455(1);
  n3857 <= tmp_ivl_11455(0);
  tmp_ivl_11455 <= LPM_d0_ivl_11459(0 + 1 downto 0);
  tmp_ivl_11461 <= z1(18);
  tmp_ivl_11462 <= new_AGEMA_signal_2999 & tmp_ivl_11461;
  LPM_q_ivl_11465 <= tmp_ivl_11467 & tmp_ivl_11462;
  tmp_ivl_11469 <= new_AGEMA_signal_3353 & n3857;
  LPM_q_ivl_11472 <= tmp_ivl_11474 & tmp_ivl_11469;
  new_AGEMA_signal_3636 <= tmp_ivl_11476(1);
  n3337 <= tmp_ivl_11476(0);
  tmp_ivl_11476 <= LPM_d0_ivl_11480(0 + 1 downto 0);
  tmp_ivl_11481 <= new_AGEMA_signal_3636 & n3337;
  LPM_q_ivl_11484 <= tmp_ivl_11486 & tmp_ivl_11481;
  tmp_ivl_11488 <= new_AGEMA_signal_2663 & n3336;
  LPM_q_ivl_11491 <= tmp_ivl_11493 & tmp_ivl_11488;
  new_AGEMA_signal_3920 <= tmp_ivl_11495(1);
  n3648 <= tmp_ivl_11495(0);
  tmp_ivl_11495 <= LPM_d0_ivl_11499(0 + 1 downto 0);
  tmp_ivl_11500 <= new_AGEMA_signal_4226 & n3338;
  LPM_q_ivl_11503 <= tmp_ivl_11505 & tmp_ivl_11500;
  tmp_ivl_11507 <= new_AGEMA_signal_3920 & n3648;
  LPM_q_ivl_11510 <= tmp_ivl_11512 & tmp_ivl_11507;
  tmp_ivl_11514 <= tmp_ivl_11518(1);
  tmp_ivl_11516 <= tmp_ivl_11518(0);
  tmp_ivl_11518 <= LPM_d0_ivl_11522(0 + 1 downto 0);
  tmp_ivl_11524 <= z1(19);
  tmp_ivl_11525 <= new_AGEMA_signal_3000 & tmp_ivl_11524;
  LPM_q_ivl_11528 <= tmp_ivl_11530 & tmp_ivl_11525;
  tmp_ivl_11533 <= state_in_s1(299);
  tmp_ivl_11535 <= state_in_s0(299);
  tmp_ivl_11536 <= tmp_ivl_11533 & tmp_ivl_11535;
  LPM_q_ivl_11539 <= tmp_ivl_11541 & tmp_ivl_11536;
  new_AGEMA_signal_3354 <= tmp_ivl_11543(1);
  n3340 <= tmp_ivl_11543(0);
  tmp_ivl_11543 <= LPM_d0_ivl_11547(0 + 1 downto 0);
  tmp_ivl_11549 <= z0(19);
  tmp_ivl_11550 <= new_AGEMA_signal_3242 & tmp_ivl_11549;
  LPM_q_ivl_11553 <= tmp_ivl_11555 & tmp_ivl_11550;
  tmp_ivl_11558 <= state_in_s1(43);
  tmp_ivl_11560 <= state_in_s0(43);
  tmp_ivl_11561 <= tmp_ivl_11558 & tmp_ivl_11560;
  LPM_q_ivl_11564 <= tmp_ivl_11566 & tmp_ivl_11561;
  new_AGEMA_signal_3355 <= tmp_ivl_11568(1);
  n3356 <= tmp_ivl_11568(0);
  tmp_ivl_11568 <= LPM_d0_ivl_11572(0 + 1 downto 0);
  tmp_ivl_11574 <= state_in_s1(107);
  tmp_ivl_11576 <= state_in_s0(107);
  tmp_ivl_11577 <= tmp_ivl_11574 & tmp_ivl_11576;
  LPM_q_ivl_11580 <= tmp_ivl_11582 & tmp_ivl_11577;
  tmp_ivl_11584 <= new_AGEMA_signal_3355 & n3356;
  LPM_q_ivl_11587 <= tmp_ivl_11589 & tmp_ivl_11584;
  new_AGEMA_signal_3637 <= tmp_ivl_11591(1);
  n3339 <= tmp_ivl_11591(0);
  tmp_ivl_11591 <= LPM_d0_ivl_11595(0 + 1 downto 0);
  tmp_ivl_11596 <= new_AGEMA_signal_3354 & n3340;
  LPM_q_ivl_11599 <= tmp_ivl_11601 & tmp_ivl_11596;
  tmp_ivl_11603 <= new_AGEMA_signal_3637 & n3339;
  LPM_q_ivl_11606 <= tmp_ivl_11608 & tmp_ivl_11603;
  new_AGEMA_signal_3921 <= tmp_ivl_11610(1);
  n3697 <= tmp_ivl_11610(0);
  tmp_ivl_11610 <= LPM_d0_ivl_11614(0 + 1 downto 0);
  tmp_ivl_11615 <= new_AGEMA_signal_3907 & n3542;
  LPM_q_ivl_11618 <= tmp_ivl_11620 & tmp_ivl_11615;
  tmp_ivl_11622 <= new_AGEMA_signal_3921 & n3697;
  LPM_q_ivl_11625 <= tmp_ivl_11627 & tmp_ivl_11622;
  new_AGEMA_signal_4227 <= tmp_ivl_11629(1);
  n3343 <= tmp_ivl_11629(0);
  tmp_ivl_11629 <= LPM_d0_ivl_11633(0 + 1 downto 0);
  tmp_ivl_11635 <= z1(16);
  tmp_ivl_11636 <= new_AGEMA_signal_2997 & tmp_ivl_11635;
  LPM_q_ivl_11639 <= tmp_ivl_11641 & tmp_ivl_11636;
  tmp_ivl_11644 <= state_in_s1(296);
  tmp_ivl_11646 <= state_in_s0(296);
  tmp_ivl_11647 <= tmp_ivl_11644 & tmp_ivl_11646;
  LPM_q_ivl_11650 <= tmp_ivl_11652 & tmp_ivl_11647;
  new_AGEMA_signal_3356 <= tmp_ivl_11654(1);
  n3342 <= tmp_ivl_11654(0);
  tmp_ivl_11654 <= LPM_d0_ivl_11658(0 + 1 downto 0);
  tmp_ivl_11660 <= z0(16);
  tmp_ivl_11661 <= new_AGEMA_signal_3250 & tmp_ivl_11660;
  LPM_q_ivl_11664 <= tmp_ivl_11666 & tmp_ivl_11661;
  tmp_ivl_11669 <= state_in_s1(40);
  tmp_ivl_11671 <= state_in_s0(40);
  tmp_ivl_11672 <= tmp_ivl_11669 & tmp_ivl_11671;
  LPM_q_ivl_11675 <= tmp_ivl_11677 & tmp_ivl_11672;
  new_AGEMA_signal_3357 <= tmp_ivl_11679(1);
  n3682 <= tmp_ivl_11679(0);
  tmp_ivl_11679 <= LPM_d0_ivl_11683(0 + 1 downto 0);
  tmp_ivl_11685 <= state_in_s1(104);
  tmp_ivl_11687 <= state_in_s0(104);
  tmp_ivl_11688 <= tmp_ivl_11685 & tmp_ivl_11687;
  LPM_q_ivl_11691 <= tmp_ivl_11693 & tmp_ivl_11688;
  tmp_ivl_11695 <= new_AGEMA_signal_3357 & n3682;
  LPM_q_ivl_11698 <= tmp_ivl_11700 & tmp_ivl_11695;
  new_AGEMA_signal_3638 <= tmp_ivl_11702(1);
  n3341 <= tmp_ivl_11702(0);
  tmp_ivl_11702 <= LPM_d0_ivl_11706(0 + 1 downto 0);
  tmp_ivl_11707 <= new_AGEMA_signal_3356 & n3342;
  LPM_q_ivl_11710 <= tmp_ivl_11712 & tmp_ivl_11707;
  tmp_ivl_11714 <= new_AGEMA_signal_3638 & n3341;
  LPM_q_ivl_11717 <= tmp_ivl_11719 & tmp_ivl_11714;
  new_AGEMA_signal_3922 <= tmp_ivl_11721(1);
  n3608 <= tmp_ivl_11721(0);
  tmp_ivl_11721 <= LPM_d0_ivl_11725(0 + 1 downto 0);
  tmp_ivl_11726 <= new_AGEMA_signal_4227 & n3343;
  LPM_q_ivl_11729 <= tmp_ivl_11731 & tmp_ivl_11726;
  tmp_ivl_11733 <= new_AGEMA_signal_3922 & n3608;
  LPM_q_ivl_11736 <= tmp_ivl_11738 & tmp_ivl_11733;
  tmp_ivl_11740 <= tmp_ivl_11744(1);
  tmp_ivl_11742 <= tmp_ivl_11744(0);
  tmp_ivl_11744 <= LPM_d0_ivl_11748(0 + 1 downto 0);
  tmp_ivl_11749 <= new_AGEMA_signal_3606 & n3457;
  LPM_q_ivl_11752 <= tmp_ivl_11754 & tmp_ivl_11749;
  tmp_ivl_11756 <= new_AGEMA_signal_3608 & n3777;
  LPM_q_ivl_11759 <= tmp_ivl_11761 & tmp_ivl_11756;
  new_AGEMA_signal_3923 <= tmp_ivl_11763(1);
  n3344 <= tmp_ivl_11763(0);
  tmp_ivl_11763 <= LPM_d0_ivl_11767(0 + 1 downto 0);
  tmp_ivl_11769 <= state_in_s1(224);
  tmp_ivl_11771 <= state_in_s0(224);
  tmp_ivl_11772 <= tmp_ivl_11769 & tmp_ivl_11771;
  LPM_q_ivl_11775 <= tmp_ivl_11777 & tmp_ivl_11772;
  tmp_ivl_11780 <= z4(24);
  tmp_ivl_11781 <= new_AGEMA_signal_3127 & tmp_ivl_11780;
  LPM_q_ivl_11784 <= tmp_ivl_11786 & tmp_ivl_11781;
  new_AGEMA_signal_3358 <= tmp_ivl_11788(1);
  n3484 <= tmp_ivl_11788(0);
  tmp_ivl_11788 <= LPM_d0_ivl_11792(0 + 1 downto 0);
  tmp_ivl_11794 <= state_in_s1(288);
  tmp_ivl_11796 <= state_in_s0(288);
  tmp_ivl_11797 <= tmp_ivl_11794 & tmp_ivl_11796;
  LPM_q_ivl_11800 <= tmp_ivl_11802 & tmp_ivl_11797;
  tmp_ivl_11804 <= new_AGEMA_signal_3358 & n3484;
  LPM_q_ivl_11807 <= tmp_ivl_11809 & tmp_ivl_11804;
  new_AGEMA_signal_3639 <= tmp_ivl_11811(1);
  n3780 <= tmp_ivl_11811(0);
  tmp_ivl_11811 <= LPM_d0_ivl_11815(0 + 1 downto 0);
  tmp_ivl_11816 <= new_AGEMA_signal_3923 & n3344;
  LPM_q_ivl_11819 <= tmp_ivl_11821 & tmp_ivl_11816;
  tmp_ivl_11823 <= new_AGEMA_signal_3639 & n3780;
  LPM_q_ivl_11826 <= tmp_ivl_11828 & tmp_ivl_11823;
  tmp_ivl_11830 <= tmp_ivl_11834(1);
  tmp_ivl_11832 <= tmp_ivl_11834(0);
  tmp_ivl_11834 <= LPM_d0_ivl_11838(0 + 1 downto 0);
  tmp_ivl_11839 <= new_AGEMA_signal_3590 & n3351;
  LPM_q_ivl_11842 <= tmp_ivl_11844 & tmp_ivl_11839;
  tmp_ivl_11846 <= new_AGEMA_signal_3629 & n3456;
  LPM_q_ivl_11849 <= tmp_ivl_11851 & tmp_ivl_11846;
  new_AGEMA_signal_3924 <= tmp_ivl_11853(1);
  n3345 <= tmp_ivl_11853(0);
  tmp_ivl_11853 <= LPM_d0_ivl_11857(0 + 1 downto 0);
  tmp_ivl_11858 <= new_AGEMA_signal_3924 & n3345;
  LPM_q_ivl_11861 <= tmp_ivl_11863 & tmp_ivl_11858;
  tmp_ivl_11865 <= new_AGEMA_signal_3639 & n3780;
  LPM_q_ivl_11868 <= tmp_ivl_11870 & tmp_ivl_11865;
  tmp_ivl_11872 <= tmp_ivl_11876(1);
  tmp_ivl_11874 <= tmp_ivl_11876(0);
  tmp_ivl_11876 <= LPM_d0_ivl_11880(0 + 1 downto 0);
  tmp_ivl_11882 <= z1(20);
  tmp_ivl_11883 <= new_AGEMA_signal_3001 & tmp_ivl_11882;
  LPM_q_ivl_11886 <= tmp_ivl_11888 & tmp_ivl_11883;
  tmp_ivl_11891 <= state_in_s1(300);
  tmp_ivl_11893 <= state_in_s0(300);
  tmp_ivl_11894 <= tmp_ivl_11891 & tmp_ivl_11893;
  LPM_q_ivl_11897 <= tmp_ivl_11899 & tmp_ivl_11894;
  new_AGEMA_signal_3359 <= tmp_ivl_11901(1);
  n3347 <= tmp_ivl_11901(0);
  tmp_ivl_11901 <= LPM_d0_ivl_11905(0 + 1 downto 0);
  tmp_ivl_11907 <= z0(20);
  tmp_ivl_11908 <= new_AGEMA_signal_3240 & tmp_ivl_11907;
  LPM_q_ivl_11911 <= tmp_ivl_11913 & tmp_ivl_11908;
  tmp_ivl_11916 <= state_in_s1(44);
  tmp_ivl_11918 <= state_in_s0(44);
  tmp_ivl_11919 <= tmp_ivl_11916 & tmp_ivl_11918;
  LPM_q_ivl_11922 <= tmp_ivl_11924 & tmp_ivl_11919;
  new_AGEMA_signal_3360 <= tmp_ivl_11926(1);
  n3440 <= tmp_ivl_11926(0);
  tmp_ivl_11926 <= LPM_d0_ivl_11930(0 + 1 downto 0);
  tmp_ivl_11932 <= state_in_s1(108);
  tmp_ivl_11934 <= state_in_s0(108);
  tmp_ivl_11935 <= tmp_ivl_11932 & tmp_ivl_11934;
  LPM_q_ivl_11938 <= tmp_ivl_11940 & tmp_ivl_11935;
  tmp_ivl_11942 <= new_AGEMA_signal_3360 & n3440;
  LPM_q_ivl_11945 <= tmp_ivl_11947 & tmp_ivl_11942;
  new_AGEMA_signal_3640 <= tmp_ivl_11949(1);
  n3346 <= tmp_ivl_11949(0);
  tmp_ivl_11949 <= LPM_d0_ivl_11953(0 + 1 downto 0);
  tmp_ivl_11954 <= new_AGEMA_signal_3359 & n3347;
  LPM_q_ivl_11957 <= tmp_ivl_11959 & tmp_ivl_11954;
  tmp_ivl_11961 <= new_AGEMA_signal_3640 & n3346;
  LPM_q_ivl_11964 <= tmp_ivl_11966 & tmp_ivl_11961;
  new_AGEMA_signal_3925 <= tmp_ivl_11968(1);
  n3796 <= tmp_ivl_11968(0);
  tmp_ivl_11968 <= LPM_d0_ivl_11972(0 + 1 downto 0);
  tmp_ivl_11973 <= new_AGEMA_signal_3910 & n3572;
  LPM_q_ivl_11976 <= tmp_ivl_11978 & tmp_ivl_11973;
  tmp_ivl_11980 <= new_AGEMA_signal_3925 & n3796;
  LPM_q_ivl_11983 <= tmp_ivl_11985 & tmp_ivl_11980;
  new_AGEMA_signal_4230 <= tmp_ivl_11987(1);
  n3350 <= tmp_ivl_11987(0);
  tmp_ivl_11987 <= LPM_d0_ivl_11991(0 + 1 downto 0);
  tmp_ivl_11993 <= z0(17);
  tmp_ivl_11994 <= new_AGEMA_signal_3248 & tmp_ivl_11993;
  LPM_q_ivl_11997 <= tmp_ivl_11999 & tmp_ivl_11994;
  tmp_ivl_12002 <= state_in_s1(41);
  tmp_ivl_12004 <= state_in_s0(41);
  tmp_ivl_12005 <= tmp_ivl_12002 & tmp_ivl_12004;
  LPM_q_ivl_12008 <= tmp_ivl_12010 & tmp_ivl_12005;
  new_AGEMA_signal_3361 <= tmp_ivl_12012(1);
  n3771 <= tmp_ivl_12012(0);
  tmp_ivl_12012 <= LPM_d0_ivl_12016(0 + 1 downto 0);
  tmp_ivl_12018 <= z1(17);
  tmp_ivl_12019 <= new_AGEMA_signal_2998 & tmp_ivl_12018;
  LPM_q_ivl_12022 <= tmp_ivl_12024 & tmp_ivl_12019;
  tmp_ivl_12026 <= new_AGEMA_signal_3361 & n3771;
  LPM_q_ivl_12029 <= tmp_ivl_12031 & tmp_ivl_12026;
  new_AGEMA_signal_3641 <= tmp_ivl_12033(1);
  n3349 <= tmp_ivl_12033(0);
  tmp_ivl_12033 <= LPM_d0_ivl_12037(0 + 1 downto 0);
  tmp_ivl_12038 <= new_AGEMA_signal_3641 & n3349;
  LPM_q_ivl_12041 <= tmp_ivl_12043 & tmp_ivl_12038;
  tmp_ivl_12045 <= new_AGEMA_signal_2665 & n3348;
  LPM_q_ivl_12048 <= tmp_ivl_12050 & tmp_ivl_12045;
  new_AGEMA_signal_3926 <= tmp_ivl_12052(1);
  n3617 <= tmp_ivl_12052(0);
  tmp_ivl_12052 <= LPM_d0_ivl_12056(0 + 1 downto 0);
  tmp_ivl_12057 <= new_AGEMA_signal_4230 & n3350;
  LPM_q_ivl_12060 <= tmp_ivl_12062 & tmp_ivl_12057;
  tmp_ivl_12064 <= new_AGEMA_signal_3926 & n3617;
  LPM_q_ivl_12067 <= tmp_ivl_12069 & tmp_ivl_12064;
  tmp_ivl_12071 <= tmp_ivl_12075(1);
  tmp_ivl_12073 <= tmp_ivl_12075(0);
  tmp_ivl_12075 <= LPM_d0_ivl_12079(0 + 1 downto 0);
  tmp_ivl_12080 <= new_AGEMA_signal_3590 & n3351;
  LPM_q_ivl_12083 <= tmp_ivl_12085 & tmp_ivl_12080;
  tmp_ivl_12087 <= new_AGEMA_signal_3616 & n3481;
  LPM_q_ivl_12090 <= tmp_ivl_12092 & tmp_ivl_12087;
  new_AGEMA_signal_3927 <= tmp_ivl_12094(1);
  n3352 <= tmp_ivl_12094(0);
  tmp_ivl_12094 <= LPM_d0_ivl_12098(0 + 1 downto 0);
  tmp_ivl_12100 <= state_in_s1(194);
  tmp_ivl_12102 <= state_in_s0(194);
  tmp_ivl_12103 <= tmp_ivl_12100 & tmp_ivl_12102;
  LPM_q_ivl_12106 <= tmp_ivl_12108 & tmp_ivl_12103;
  tmp_ivl_12111 <= z4(58);
  tmp_ivl_12112 <= new_AGEMA_signal_3164 & tmp_ivl_12111;
  LPM_q_ivl_12115 <= tmp_ivl_12117 & tmp_ivl_12112;
  new_AGEMA_signal_3362 <= tmp_ivl_12119(1);
  n3406 <= tmp_ivl_12119(0);
  tmp_ivl_12119 <= LPM_d0_ivl_12123(0 + 1 downto 0);
  tmp_ivl_12125 <= state_in_s1(258);
  tmp_ivl_12127 <= state_in_s0(258);
  tmp_ivl_12128 <= tmp_ivl_12125 & tmp_ivl_12127;
  LPM_q_ivl_12131 <= tmp_ivl_12133 & tmp_ivl_12128;
  tmp_ivl_12135 <= new_AGEMA_signal_3362 & n3406;
  LPM_q_ivl_12138 <= tmp_ivl_12140 & tmp_ivl_12135;
  new_AGEMA_signal_3642 <= tmp_ivl_12142(1);
  n3832 <= tmp_ivl_12142(0);
  tmp_ivl_12142 <= LPM_d0_ivl_12146(0 + 1 downto 0);
  tmp_ivl_12147 <= new_AGEMA_signal_3927 & n3352;
  LPM_q_ivl_12150 <= tmp_ivl_12152 & tmp_ivl_12147;
  tmp_ivl_12154 <= new_AGEMA_signal_3642 & n3832;
  LPM_q_ivl_12157 <= tmp_ivl_12159 & tmp_ivl_12154;
  tmp_ivl_12161 <= tmp_ivl_12165(1);
  tmp_ivl_12163 <= tmp_ivl_12165(0);
  tmp_ivl_12165 <= LPM_d0_ivl_12169(0 + 1 downto 0);
  tmp_ivl_12171 <= z0(38);
  tmp_ivl_12172 <= new_AGEMA_signal_3264 & tmp_ivl_12171;
  LPM_q_ivl_12175 <= tmp_ivl_12177 & tmp_ivl_12172;
  tmp_ivl_12180 <= state_in_s1(30);
  tmp_ivl_12182 <= state_in_s0(30);
  tmp_ivl_12183 <= tmp_ivl_12180 & tmp_ivl_12182;
  LPM_q_ivl_12186 <= tmp_ivl_12188 & tmp_ivl_12183;
  new_AGEMA_signal_3363 <= tmp_ivl_12190(1);
  n3409 <= tmp_ivl_12190(0);
  tmp_ivl_12190 <= LPM_d0_ivl_12194(0 + 1 downto 0);
  tmp_ivl_12195 <= new_AGEMA_signal_3363 & n3409;
  LPM_q_ivl_12198 <= tmp_ivl_12200 & tmp_ivl_12195;
  tmp_ivl_12202 <= new_AGEMA_signal_3342 & n3353;
  LPM_q_ivl_12205 <= tmp_ivl_12207 & tmp_ivl_12202;
  new_AGEMA_signal_3643 <= tmp_ivl_12209(1);
  n3709 <= tmp_ivl_12209(0);
  tmp_ivl_12209 <= LPM_d0_ivl_12213(0 + 1 downto 0);
  tmp_ivl_12215 <= z0(47);
  tmp_ivl_12216 <= new_AGEMA_signal_3239 & tmp_ivl_12215;
  LPM_q_ivl_12219 <= tmp_ivl_12221 & tmp_ivl_12216;
  tmp_ivl_12224 <= state_in_s1(23);
  tmp_ivl_12226 <= state_in_s0(23);
  tmp_ivl_12227 <= tmp_ivl_12224 & tmp_ivl_12226;
  LPM_q_ivl_12230 <= tmp_ivl_12232 & tmp_ivl_12227;
  new_AGEMA_signal_3364 <= tmp_ivl_12234(1);
  n3369 <= tmp_ivl_12234(0);
  tmp_ivl_12234 <= LPM_d0_ivl_12238(0 + 1 downto 0);
  tmp_ivl_12239 <= new_AGEMA_signal_3364 & n3369;
  LPM_q_ivl_12242 <= tmp_ivl_12244 & tmp_ivl_12239;
  tmp_ivl_12246 <= new_AGEMA_signal_3318 & n3354;
  LPM_q_ivl_12249 <= tmp_ivl_12251 & tmp_ivl_12246;
  new_AGEMA_signal_3644 <= tmp_ivl_12253(1);
  n3705 <= tmp_ivl_12253(0);
  tmp_ivl_12253 <= LPM_d0_ivl_12257(0 + 1 downto 0);
  tmp_ivl_12258 <= new_AGEMA_signal_3643 & n3709;
  LPM_q_ivl_12261 <= tmp_ivl_12263 & tmp_ivl_12258;
  tmp_ivl_12265 <= new_AGEMA_signal_3644 & n3705;
  LPM_q_ivl_12268 <= tmp_ivl_12270 & tmp_ivl_12265;
  new_AGEMA_signal_3928 <= tmp_ivl_12272(1);
  n3357 <= tmp_ivl_12272(0);
  tmp_ivl_12272 <= LPM_d0_ivl_12276(0 + 1 downto 0);
  tmp_ivl_12277 <= new_AGEMA_signal_3355 & n3356;
  LPM_q_ivl_12280 <= tmp_ivl_12282 & tmp_ivl_12277;
  tmp_ivl_12284 <= new_AGEMA_signal_3310 & n3355;
  LPM_q_ivl_12287 <= tmp_ivl_12289 & tmp_ivl_12284;
  new_AGEMA_signal_3645 <= tmp_ivl_12291(1);
  n3637 <= tmp_ivl_12291(0);
  tmp_ivl_12291 <= LPM_d0_ivl_12295(0 + 1 downto 0);
  tmp_ivl_12296 <= new_AGEMA_signal_3928 & n3357;
  LPM_q_ivl_12299 <= tmp_ivl_12301 & tmp_ivl_12296;
  tmp_ivl_12303 <= new_AGEMA_signal_3645 & n3637;
  LPM_q_ivl_12306 <= tmp_ivl_12308 & tmp_ivl_12303;
  tmp_ivl_12310 <= tmp_ivl_12314(1);
  tmp_ivl_12312 <= tmp_ivl_12314(0);
  tmp_ivl_12314 <= LPM_d0_ivl_12318(0 + 1 downto 0);
  tmp_ivl_12320 <= state_in_s1(225);
  tmp_ivl_12322 <= state_in_s0(225);
  tmp_ivl_12323 <= tmp_ivl_12320 & tmp_ivl_12322;
  LPM_q_ivl_12326 <= tmp_ivl_12328 & tmp_ivl_12323;
  tmp_ivl_12331 <= z4(25);
  tmp_ivl_12332 <= new_AGEMA_signal_3128 & tmp_ivl_12331;
  LPM_q_ivl_12335 <= tmp_ivl_12337 & tmp_ivl_12332;
  new_AGEMA_signal_3365 <= tmp_ivl_12339(1);
  n3683 <= tmp_ivl_12339(0);
  tmp_ivl_12339 <= LPM_d0_ivl_12343(0 + 1 downto 0);
  tmp_ivl_12345 <= state_in_s1(289);
  tmp_ivl_12347 <= state_in_s0(289);
  tmp_ivl_12348 <= tmp_ivl_12345 & tmp_ivl_12347;
  LPM_q_ivl_12351 <= tmp_ivl_12353 & tmp_ivl_12348;
  tmp_ivl_12355 <= new_AGEMA_signal_3365 & n3683;
  LPM_q_ivl_12358 <= tmp_ivl_12360 & tmp_ivl_12355;
  new_AGEMA_signal_3646 <= tmp_ivl_12362(1);
  n3870 <= tmp_ivl_12362(0);
  tmp_ivl_12362 <= LPM_d0_ivl_12366(0 + 1 downto 0);
  tmp_ivl_12367 <= new_AGEMA_signal_3621 & n3510;
  LPM_q_ivl_12370 <= tmp_ivl_12372 & tmp_ivl_12367;
  tmp_ivl_12374 <= new_AGEMA_signal_3646 & n3870;
  LPM_q_ivl_12377 <= tmp_ivl_12379 & tmp_ivl_12374;
  new_AGEMA_signal_3929 <= tmp_ivl_12381(1);
  n3358 <= tmp_ivl_12381(0);
  tmp_ivl_12381 <= LPM_d0_ivl_12385(0 + 1 downto 0);
  tmp_ivl_12387 <= state_in_s1(200);
  tmp_ivl_12389 <= state_in_s0(200);
  tmp_ivl_12390 <= tmp_ivl_12387 & tmp_ivl_12389;
  LPM_q_ivl_12393 <= tmp_ivl_12395 & tmp_ivl_12390;
  tmp_ivl_12398 <= z4(48);
  tmp_ivl_12399 <= new_AGEMA_signal_3153 & tmp_ivl_12398;
  LPM_q_ivl_12402 <= tmp_ivl_12404 & tmp_ivl_12399;
  new_AGEMA_signal_3366 <= tmp_ivl_12406(1);
  n3527 <= tmp_ivl_12406(0);
  tmp_ivl_12406 <= LPM_d0_ivl_12410(0 + 1 downto 0);
  tmp_ivl_12412 <= state_in_s1(264);
  tmp_ivl_12414 <= state_in_s0(264);
  tmp_ivl_12415 <= tmp_ivl_12412 & tmp_ivl_12414;
  LPM_q_ivl_12418 <= tmp_ivl_12420 & tmp_ivl_12415;
  tmp_ivl_12422 <= new_AGEMA_signal_3366 & n3527;
  LPM_q_ivl_12425 <= tmp_ivl_12427 & tmp_ivl_12422;
  new_AGEMA_signal_3647 <= tmp_ivl_12429(1);
  n3866 <= tmp_ivl_12429(0);
  tmp_ivl_12429 <= LPM_d0_ivl_12433(0 + 1 downto 0);
  tmp_ivl_12434 <= new_AGEMA_signal_3929 & n3358;
  LPM_q_ivl_12437 <= tmp_ivl_12439 & tmp_ivl_12434;
  tmp_ivl_12441 <= new_AGEMA_signal_3647 & n3866;
  LPM_q_ivl_12444 <= tmp_ivl_12446 & tmp_ivl_12441;
  tmp_ivl_12448 <= tmp_ivl_12452(1);
  tmp_ivl_12450 <= tmp_ivl_12452(0);
  tmp_ivl_12452 <= LPM_d0_ivl_12456(0 + 1 downto 0);
  tmp_ivl_12457 <= new_AGEMA_signal_3593 & n3360;
  LPM_q_ivl_12460 <= tmp_ivl_12462 & tmp_ivl_12457;
  tmp_ivl_12464 <= new_AGEMA_signal_3611 & n3511;
  LPM_q_ivl_12467 <= tmp_ivl_12469 & tmp_ivl_12464;
  new_AGEMA_signal_3930 <= tmp_ivl_12471(1);
  n3359 <= tmp_ivl_12471(0);
  tmp_ivl_12471 <= LPM_d0_ivl_12475(0 + 1 downto 0);
  tmp_ivl_12476 <= new_AGEMA_signal_3930 & n3359;
  LPM_q_ivl_12479 <= tmp_ivl_12481 & tmp_ivl_12476;
  tmp_ivl_12483 <= new_AGEMA_signal_3646 & n3870;
  LPM_q_ivl_12486 <= tmp_ivl_12488 & tmp_ivl_12483;
  tmp_ivl_12490 <= tmp_ivl_12494(1);
  tmp_ivl_12492 <= tmp_ivl_12494(0);
  tmp_ivl_12494 <= LPM_d0_ivl_12498(0 + 1 downto 0);
  tmp_ivl_12499 <= new_AGEMA_signal_3593 & n3360;
  LPM_q_ivl_12502 <= tmp_ivl_12504 & tmp_ivl_12499;
  tmp_ivl_12506 <= new_AGEMA_signal_3617 & n3538;
  LPM_q_ivl_12509 <= tmp_ivl_12511 & tmp_ivl_12506;
  new_AGEMA_signal_3931 <= tmp_ivl_12513(1);
  n3361 <= tmp_ivl_12513(0);
  tmp_ivl_12513 <= LPM_d0_ivl_12517(0 + 1 downto 0);
  tmp_ivl_12519 <= state_in_s1(195);
  tmp_ivl_12521 <= state_in_s0(195);
  tmp_ivl_12522 <= tmp_ivl_12519 & tmp_ivl_12521;
  LPM_q_ivl_12525 <= tmp_ivl_12527 & tmp_ivl_12522;
  tmp_ivl_12530 <= z4(59);
  tmp_ivl_12531 <= new_AGEMA_signal_3165 & tmp_ivl_12530;
  LPM_q_ivl_12534 <= tmp_ivl_12536 & tmp_ivl_12531;
  new_AGEMA_signal_3367 <= tmp_ivl_12538(1);
  n3596 <= tmp_ivl_12538(0);
  tmp_ivl_12538 <= LPM_d0_ivl_12542(0 + 1 downto 0);
  tmp_ivl_12544 <= state_in_s1(259);
  tmp_ivl_12546 <= state_in_s0(259);
  tmp_ivl_12547 <= tmp_ivl_12544 & tmp_ivl_12546;
  LPM_q_ivl_12550 <= tmp_ivl_12552 & tmp_ivl_12547;
  tmp_ivl_12554 <= new_AGEMA_signal_3367 & n3596;
  LPM_q_ivl_12557 <= tmp_ivl_12559 & tmp_ivl_12554;
  new_AGEMA_signal_3648 <= tmp_ivl_12561(1);
  n3922 <= tmp_ivl_12561(0);
  tmp_ivl_12561 <= LPM_d0_ivl_12565(0 + 1 downto 0);
  tmp_ivl_12566 <= new_AGEMA_signal_3931 & n3361;
  LPM_q_ivl_12569 <= tmp_ivl_12571 & tmp_ivl_12566;
  tmp_ivl_12573 <= new_AGEMA_signal_3648 & n3922;
  LPM_q_ivl_12576 <= tmp_ivl_12578 & tmp_ivl_12573;
  tmp_ivl_12580 <= tmp_ivl_12584(1);
  tmp_ivl_12582 <= tmp_ivl_12584(0);
  tmp_ivl_12584 <= LPM_d0_ivl_12588(0 + 1 downto 0);
  tmp_ivl_12590 <= z1(8);
  tmp_ivl_12591 <= new_AGEMA_signal_3045 & tmp_ivl_12590;
  LPM_q_ivl_12594 <= tmp_ivl_12596 & tmp_ivl_12591;
  tmp_ivl_12599 <= state_in_s1(304);
  tmp_ivl_12601 <= state_in_s0(304);
  tmp_ivl_12602 <= tmp_ivl_12599 & tmp_ivl_12601;
  LPM_q_ivl_12605 <= tmp_ivl_12607 & tmp_ivl_12602;
  new_AGEMA_signal_3368 <= tmp_ivl_12609(1);
  n3363 <= tmp_ivl_12609(0);
  tmp_ivl_12609 <= LPM_d0_ivl_12613(0 + 1 downto 0);
  tmp_ivl_12615 <= z0(8);
  tmp_ivl_12616 <= new_AGEMA_signal_3235 & tmp_ivl_12615;
  LPM_q_ivl_12619 <= tmp_ivl_12621 & tmp_ivl_12616;
  tmp_ivl_12624 <= state_in_s1(48);
  tmp_ivl_12626 <= state_in_s0(48);
  tmp_ivl_12627 <= tmp_ivl_12624 & tmp_ivl_12626;
  LPM_q_ivl_12630 <= tmp_ivl_12632 & tmp_ivl_12627;
  new_AGEMA_signal_3369 <= tmp_ivl_12634(1);
  n3420 <= tmp_ivl_12634(0);
  tmp_ivl_12634 <= LPM_d0_ivl_12638(0 + 1 downto 0);
  tmp_ivl_12640 <= state_in_s1(112);
  tmp_ivl_12642 <= state_in_s0(112);
  tmp_ivl_12643 <= tmp_ivl_12640 & tmp_ivl_12642;
  LPM_q_ivl_12646 <= tmp_ivl_12648 & tmp_ivl_12643;
  tmp_ivl_12650 <= new_AGEMA_signal_3369 & n3420;
  LPM_q_ivl_12653 <= tmp_ivl_12655 & tmp_ivl_12650;
  new_AGEMA_signal_3649 <= tmp_ivl_12657(1);
  n3362 <= tmp_ivl_12657(0);
  tmp_ivl_12657 <= LPM_d0_ivl_12661(0 + 1 downto 0);
  tmp_ivl_12662 <= new_AGEMA_signal_3368 & n3363;
  LPM_q_ivl_12665 <= tmp_ivl_12667 & tmp_ivl_12662;
  tmp_ivl_12669 <= new_AGEMA_signal_3649 & n3362;
  LPM_q_ivl_12672 <= tmp_ivl_12674 & tmp_ivl_12669;
  new_AGEMA_signal_3932 <= tmp_ivl_12676(1);
  n3751 <= tmp_ivl_12676(0);
  tmp_ivl_12676 <= LPM_d0_ivl_12680(0 + 1 downto 0);
  tmp_ivl_12681 <= new_AGEMA_signal_3908 & n3447;
  LPM_q_ivl_12684 <= tmp_ivl_12686 & tmp_ivl_12681;
  tmp_ivl_12688 <= new_AGEMA_signal_3932 & n3751;
  LPM_q_ivl_12691 <= tmp_ivl_12693 & tmp_ivl_12688;
  new_AGEMA_signal_4236 <= tmp_ivl_12695(1);
  n3366 <= tmp_ivl_12695(0);
  tmp_ivl_12695 <= LPM_d0_ivl_12699(0 + 1 downto 0);
  tmp_ivl_12701 <= z1(30);
  tmp_ivl_12702 <= new_AGEMA_signal_3011 & tmp_ivl_12701;
  LPM_q_ivl_12705 <= tmp_ivl_12707 & tmp_ivl_12702;
  tmp_ivl_12710 <= state_in_s1(294);
  tmp_ivl_12712 <= state_in_s0(294);
  tmp_ivl_12713 <= tmp_ivl_12710 & tmp_ivl_12712;
  LPM_q_ivl_12716 <= tmp_ivl_12718 & tmp_ivl_12713;
  new_AGEMA_signal_3370 <= tmp_ivl_12720(1);
  n3365 <= tmp_ivl_12720(0);
  tmp_ivl_12720 <= LPM_d0_ivl_12724(0 + 1 downto 0);
  tmp_ivl_12726 <= z0(30);
  tmp_ivl_12727 <= new_AGEMA_signal_3256 & tmp_ivl_12726;
  LPM_q_ivl_12730 <= tmp_ivl_12732 & tmp_ivl_12727;
  tmp_ivl_12735 <= state_in_s1(38);
  tmp_ivl_12737 <= state_in_s0(38);
  tmp_ivl_12738 <= tmp_ivl_12735 & tmp_ivl_12737;
  LPM_q_ivl_12741 <= tmp_ivl_12743 & tmp_ivl_12738;
  new_AGEMA_signal_3371 <= tmp_ivl_12745(1);
  n3622 <= tmp_ivl_12745(0);
  tmp_ivl_12745 <= LPM_d0_ivl_12749(0 + 1 downto 0);
  tmp_ivl_12751 <= state_in_s1(102);
  tmp_ivl_12753 <= state_in_s0(102);
  tmp_ivl_12754 <= tmp_ivl_12751 & tmp_ivl_12753;
  LPM_q_ivl_12757 <= tmp_ivl_12759 & tmp_ivl_12754;
  tmp_ivl_12761 <= new_AGEMA_signal_3371 & n3622;
  LPM_q_ivl_12764 <= tmp_ivl_12766 & tmp_ivl_12761;
  new_AGEMA_signal_3650 <= tmp_ivl_12768(1);
  n3364 <= tmp_ivl_12768(0);
  tmp_ivl_12768 <= LPM_d0_ivl_12772(0 + 1 downto 0);
  tmp_ivl_12773 <= new_AGEMA_signal_3370 & n3365;
  LPM_q_ivl_12776 <= tmp_ivl_12778 & tmp_ivl_12773;
  tmp_ivl_12780 <= new_AGEMA_signal_3650 & n3364;
  LPM_q_ivl_12783 <= tmp_ivl_12785 & tmp_ivl_12780;
  new_AGEMA_signal_3933 <= tmp_ivl_12787(1);
  n3745 <= tmp_ivl_12787(0);
  tmp_ivl_12787 <= LPM_d0_ivl_12791(0 + 1 downto 0);
  tmp_ivl_12792 <= new_AGEMA_signal_4236 & n3366;
  LPM_q_ivl_12795 <= tmp_ivl_12797 & tmp_ivl_12792;
  tmp_ivl_12799 <= new_AGEMA_signal_3933 & n3745;
  LPM_q_ivl_12802 <= tmp_ivl_12804 & tmp_ivl_12799;
  tmp_ivl_12806 <= tmp_ivl_12810(1);
  tmp_ivl_12808 <= tmp_ivl_12810(0);
  tmp_ivl_12810 <= LPM_d0_ivl_12814(0 + 1 downto 0);
  tmp_ivl_12816 <= z0(25);
  tmp_ivl_12817 <= new_AGEMA_signal_3260 & tmp_ivl_12816;
  LPM_q_ivl_12820 <= tmp_ivl_12822 & tmp_ivl_12817;
  tmp_ivl_12825 <= state_in_s1(33);
  tmp_ivl_12827 <= state_in_s0(33);
  tmp_ivl_12828 <= tmp_ivl_12825 & tmp_ivl_12827;
  LPM_q_ivl_12831 <= tmp_ivl_12833 & tmp_ivl_12828;
  new_AGEMA_signal_3372 <= tmp_ivl_12835(1);
  n3684 <= tmp_ivl_12835(0);
  tmp_ivl_12835 <= LPM_d0_ivl_12839(0 + 1 downto 0);
  tmp_ivl_12841 <= z1(25);
  tmp_ivl_12842 <= new_AGEMA_signal_3006 & tmp_ivl_12841;
  LPM_q_ivl_12845 <= tmp_ivl_12847 & tmp_ivl_12842;
  tmp_ivl_12849 <= new_AGEMA_signal_3372 & n3684;
  LPM_q_ivl_12852 <= tmp_ivl_12854 & tmp_ivl_12849;
  new_AGEMA_signal_3651 <= tmp_ivl_12856(1);
  n3368 <= tmp_ivl_12856(0);
  tmp_ivl_12856 <= LPM_d0_ivl_12860(0 + 1 downto 0);
  tmp_ivl_12861 <= new_AGEMA_signal_3651 & n3368;
  LPM_q_ivl_12864 <= tmp_ivl_12866 & tmp_ivl_12861;
  tmp_ivl_12868 <= new_AGEMA_signal_2667 & n3367;
  LPM_q_ivl_12871 <= tmp_ivl_12873 & tmp_ivl_12868;
  new_AGEMA_signal_3934 <= tmp_ivl_12875(1);
  n3810 <= tmp_ivl_12875(0);
  tmp_ivl_12875 <= LPM_d0_ivl_12879(0 + 1 downto 0);
  tmp_ivl_12881 <= z1(47);
  tmp_ivl_12882 <= new_AGEMA_signal_3028 & tmp_ivl_12881;
  LPM_q_ivl_12885 <= tmp_ivl_12887 & tmp_ivl_12882;
  tmp_ivl_12889 <= new_AGEMA_signal_3364 & n3369;
  LPM_q_ivl_12892 <= tmp_ivl_12894 & tmp_ivl_12889;
  new_AGEMA_signal_3652 <= tmp_ivl_12896(1);
  n3371 <= tmp_ivl_12896(0);
  tmp_ivl_12896 <= LPM_d0_ivl_12900(0 + 1 downto 0);
  tmp_ivl_12901 <= new_AGEMA_signal_3652 & n3371;
  LPM_q_ivl_12904 <= tmp_ivl_12906 & tmp_ivl_12901;
  tmp_ivl_12908 <= new_AGEMA_signal_2669 & n3370;
  LPM_q_ivl_12911 <= tmp_ivl_12913 & tmp_ivl_12908;
  new_AGEMA_signal_3935 <= tmp_ivl_12915(1);
  n3750 <= tmp_ivl_12915(0);
  tmp_ivl_12915 <= LPM_d0_ivl_12919(0 + 1 downto 0);
  tmp_ivl_12920 <= new_AGEMA_signal_3934 & n3810;
  LPM_q_ivl_12923 <= tmp_ivl_12925 & tmp_ivl_12920;
  tmp_ivl_12927 <= new_AGEMA_signal_3935 & n3750;
  LPM_q_ivl_12930 <= tmp_ivl_12932 & tmp_ivl_12927;
  new_AGEMA_signal_4237 <= tmp_ivl_12934(1);
  n3374 <= tmp_ivl_12934(0);
  tmp_ivl_12934 <= LPM_d0_ivl_12938(0 + 1 downto 0);
  tmp_ivl_12940 <= z1(50);
  tmp_ivl_12941 <= new_AGEMA_signal_3031 & tmp_ivl_12940;
  LPM_q_ivl_12944 <= tmp_ivl_12946 & tmp_ivl_12941;
  tmp_ivl_12949 <= state_in_s1(266);
  tmp_ivl_12951 <= state_in_s0(266);
  tmp_ivl_12952 <= tmp_ivl_12949 & tmp_ivl_12951;
  LPM_q_ivl_12955 <= tmp_ivl_12957 & tmp_ivl_12952;
  new_AGEMA_signal_3373 <= tmp_ivl_12959(1);
  n3373 <= tmp_ivl_12959(0);
  tmp_ivl_12959 <= LPM_d0_ivl_12963(0 + 1 downto 0);
  tmp_ivl_12965 <= z0(50);
  tmp_ivl_12966 <= new_AGEMA_signal_3236 & tmp_ivl_12965;
  LPM_q_ivl_12969 <= tmp_ivl_12971 & tmp_ivl_12966;
  tmp_ivl_12974 <= state_in_s1(10);
  tmp_ivl_12976 <= state_in_s0(10);
  tmp_ivl_12977 <= tmp_ivl_12974 & tmp_ivl_12976;
  LPM_q_ivl_12980 <= tmp_ivl_12982 & tmp_ivl_12977;
  new_AGEMA_signal_3374 <= tmp_ivl_12984(1);
  n3722 <= tmp_ivl_12984(0);
  tmp_ivl_12984 <= LPM_d0_ivl_12988(0 + 1 downto 0);
  tmp_ivl_12990 <= state_in_s1(74);
  tmp_ivl_12992 <= state_in_s0(74);
  tmp_ivl_12993 <= tmp_ivl_12990 & tmp_ivl_12992;
  LPM_q_ivl_12996 <= tmp_ivl_12998 & tmp_ivl_12993;
  tmp_ivl_13000 <= new_AGEMA_signal_3374 & n3722;
  LPM_q_ivl_13003 <= tmp_ivl_13005 & tmp_ivl_13000;
  new_AGEMA_signal_3653 <= tmp_ivl_13007(1);
  n3372 <= tmp_ivl_13007(0);
  tmp_ivl_13007 <= LPM_d0_ivl_13011(0 + 1 downto 0);
  tmp_ivl_13012 <= new_AGEMA_signal_3373 & n3373;
  LPM_q_ivl_13015 <= tmp_ivl_13017 & tmp_ivl_13012;
  tmp_ivl_13019 <= new_AGEMA_signal_3653 & n3372;
  LPM_q_ivl_13022 <= tmp_ivl_13024 & tmp_ivl_13019;
  new_AGEMA_signal_3936 <= tmp_ivl_13026(1);
  n3468 <= tmp_ivl_13026(0);
  tmp_ivl_13026 <= LPM_d0_ivl_13030(0 + 1 downto 0);
  tmp_ivl_13031 <= new_AGEMA_signal_4237 & n3374;
  LPM_q_ivl_13034 <= tmp_ivl_13036 & tmp_ivl_13031;
  tmp_ivl_13038 <= new_AGEMA_signal_3936 & n3468;
  LPM_q_ivl_13041 <= tmp_ivl_13043 & tmp_ivl_13038;
  tmp_ivl_13045 <= tmp_ivl_13049(1);
  tmp_ivl_13047 <= tmp_ivl_13049(0);
  tmp_ivl_13049 <= LPM_d0_ivl_13053(0 + 1 downto 0);
  tmp_ivl_13054 <= new_AGEMA_signal_3596 & n3391;
  LPM_q_ivl_13057 <= tmp_ivl_13059 & tmp_ivl_13054;
  tmp_ivl_13061 <= new_AGEMA_signal_3613 & n3559;
  LPM_q_ivl_13064 <= tmp_ivl_13066 & tmp_ivl_13061;
  new_AGEMA_signal_3937 <= tmp_ivl_13068(1);
  n3375 <= tmp_ivl_13068(0);
  tmp_ivl_13068 <= LPM_d0_ivl_13072(0 + 1 downto 0);
  tmp_ivl_13074 <= state_in_s1(226);
  tmp_ivl_13076 <= state_in_s0(226);
  tmp_ivl_13077 <= tmp_ivl_13074 & tmp_ivl_13076;
  LPM_q_ivl_13080 <= tmp_ivl_13082 & tmp_ivl_13077;
  tmp_ivl_13085 <= z4(26);
  tmp_ivl_13086 <= new_AGEMA_signal_3129 & tmp_ivl_13085;
  LPM_q_ivl_13089 <= tmp_ivl_13091 & tmp_ivl_13086;
  new_AGEMA_signal_3375 <= tmp_ivl_13093(1);
  n3769 <= tmp_ivl_13093(0);
  tmp_ivl_13093 <= LPM_d0_ivl_13097(0 + 1 downto 0);
  tmp_ivl_13099 <= state_in_s1(290);
  tmp_ivl_13101 <= state_in_s0(290);
  tmp_ivl_13102 <= tmp_ivl_13099 & tmp_ivl_13101;
  LPM_q_ivl_13105 <= tmp_ivl_13107 & tmp_ivl_13102;
  tmp_ivl_13109 <= new_AGEMA_signal_3375 & n3769;
  LPM_q_ivl_13112 <= tmp_ivl_13114 & tmp_ivl_13109;
  new_AGEMA_signal_3654 <= tmp_ivl_13116(1);
  n3656 <= tmp_ivl_13116(0);
  tmp_ivl_13116 <= LPM_d0_ivl_13120(0 + 1 downto 0);
  tmp_ivl_13121 <= new_AGEMA_signal_3937 & n3375;
  LPM_q_ivl_13124 <= tmp_ivl_13126 & tmp_ivl_13121;
  tmp_ivl_13128 <= new_AGEMA_signal_3654 & n3656;
  LPM_q_ivl_13131 <= tmp_ivl_13133 & tmp_ivl_13128;
  tmp_ivl_13135 <= tmp_ivl_13139(1);
  tmp_ivl_13137 <= tmp_ivl_13139(0);
  tmp_ivl_13139 <= LPM_d0_ivl_13143(0 + 1 downto 0);
  tmp_ivl_13144 <= new_AGEMA_signal_3614 & n3867;
  LPM_q_ivl_13147 <= tmp_ivl_13149 & tmp_ivl_13144;
  tmp_ivl_13151 <= new_AGEMA_signal_3631 & n3631;
  LPM_q_ivl_13154 <= tmp_ivl_13156 & tmp_ivl_13151;
  new_AGEMA_signal_3938 <= tmp_ivl_13158(1);
  n3376 <= tmp_ivl_13158(0);
  tmp_ivl_13158 <= LPM_d0_ivl_13162(0 + 1 downto 0);
  tmp_ivl_13164 <= state_in_s1(255);
  tmp_ivl_13166 <= state_in_s0(255);
  tmp_ivl_13167 <= tmp_ivl_13164 & tmp_ivl_13166;
  LPM_q_ivl_13170 <= tmp_ivl_13172 & tmp_ivl_13167;
  tmp_ivl_13175 <= z4(7);
  tmp_ivl_13176 <= new_AGEMA_signal_3172 & tmp_ivl_13175;
  LPM_q_ivl_13179 <= tmp_ivl_13181 & tmp_ivl_13176;
  new_AGEMA_signal_3376 <= tmp_ivl_13183(1);
  n3873 <= tmp_ivl_13183(0);
  tmp_ivl_13183 <= LPM_d0_ivl_13187(0 + 1 downto 0);
  tmp_ivl_13189 <= state_in_s1(319);
  tmp_ivl_13191 <= state_in_s0(319);
  tmp_ivl_13192 <= tmp_ivl_13189 & tmp_ivl_13191;
  LPM_q_ivl_13195 <= tmp_ivl_13197 & tmp_ivl_13192;
  tmp_ivl_13199 <= new_AGEMA_signal_3376 & n3873;
  LPM_q_ivl_13202 <= tmp_ivl_13204 & tmp_ivl_13199;
  new_AGEMA_signal_3655 <= tmp_ivl_13206(1);
  n3628 <= tmp_ivl_13206(0);
  tmp_ivl_13206 <= LPM_d0_ivl_13210(0 + 1 downto 0);
  tmp_ivl_13211 <= new_AGEMA_signal_3938 & n3376;
  LPM_q_ivl_13214 <= tmp_ivl_13216 & tmp_ivl_13211;
  tmp_ivl_13218 <= new_AGEMA_signal_3655 & n3628;
  LPM_q_ivl_13221 <= tmp_ivl_13223 & tmp_ivl_13218;
  tmp_ivl_13225 <= tmp_ivl_13229(1);
  tmp_ivl_13227 <= tmp_ivl_13229(0);
  tmp_ivl_13229 <= LPM_d0_ivl_13233(0 + 1 downto 0);
  tmp_ivl_13234 <= new_AGEMA_signal_3619 & n3377;
  LPM_q_ivl_13237 <= tmp_ivl_13239 & tmp_ivl_13234;
  tmp_ivl_13241 <= new_AGEMA_signal_3647 & n3866;
  LPM_q_ivl_13244 <= tmp_ivl_13246 & tmp_ivl_13241;
  new_AGEMA_signal_3939 <= tmp_ivl_13248(1);
  n3378 <= tmp_ivl_13248(0);
  tmp_ivl_13248 <= LPM_d0_ivl_13252(0 + 1 downto 0);
  tmp_ivl_13253 <= new_AGEMA_signal_3939 & n3378;
  LPM_q_ivl_13256 <= tmp_ivl_13258 & tmp_ivl_13253;
  tmp_ivl_13260 <= new_AGEMA_signal_3655 & n3628;
  LPM_q_ivl_13263 <= tmp_ivl_13265 & tmp_ivl_13260;
  tmp_ivl_13267 <= tmp_ivl_13271(1);
  tmp_ivl_13269 <= tmp_ivl_13271(0);
  tmp_ivl_13271 <= LPM_d0_ivl_13275(0 + 1 downto 0);
  tmp_ivl_13277 <= z1(9);
  tmp_ivl_13278 <= new_AGEMA_signal_3046 & tmp_ivl_13277;
  LPM_q_ivl_13281 <= tmp_ivl_13283 & tmp_ivl_13278;
  tmp_ivl_13286 <= state_in_s1(305);
  tmp_ivl_13288 <= state_in_s0(305);
  tmp_ivl_13289 <= tmp_ivl_13286 & tmp_ivl_13288;
  LPM_q_ivl_13292 <= tmp_ivl_13294 & tmp_ivl_13289;
  new_AGEMA_signal_3377 <= tmp_ivl_13296(1);
  n3380 <= tmp_ivl_13296(0);
  tmp_ivl_13296 <= LPM_d0_ivl_13300(0 + 1 downto 0);
  tmp_ivl_13302 <= z0(9);
  tmp_ivl_13303 <= new_AGEMA_signal_3233 & tmp_ivl_13302;
  LPM_q_ivl_13306 <= tmp_ivl_13308 & tmp_ivl_13303;
  tmp_ivl_13311 <= state_in_s1(49);
  tmp_ivl_13313 <= state_in_s0(49);
  tmp_ivl_13314 <= tmp_ivl_13311 & tmp_ivl_13313;
  LPM_q_ivl_13317 <= tmp_ivl_13319 & tmp_ivl_13314;
  new_AGEMA_signal_3378 <= tmp_ivl_13321(1);
  n3479 <= tmp_ivl_13321(0);
  tmp_ivl_13321 <= LPM_d0_ivl_13325(0 + 1 downto 0);
  tmp_ivl_13327 <= state_in_s1(113);
  tmp_ivl_13329 <= state_in_s0(113);
  tmp_ivl_13330 <= tmp_ivl_13327 & tmp_ivl_13329;
  LPM_q_ivl_13333 <= tmp_ivl_13335 & tmp_ivl_13330;
  tmp_ivl_13337 <= new_AGEMA_signal_3378 & n3479;
  LPM_q_ivl_13340 <= tmp_ivl_13342 & tmp_ivl_13337;
  new_AGEMA_signal_3656 <= tmp_ivl_13344(1);
  n3379 <= tmp_ivl_13344(0);
  tmp_ivl_13344 <= LPM_d0_ivl_13348(0 + 1 downto 0);
  tmp_ivl_13349 <= new_AGEMA_signal_3377 & n3380;
  LPM_q_ivl_13352 <= tmp_ivl_13354 & tmp_ivl_13349;
  tmp_ivl_13356 <= new_AGEMA_signal_3656 & n3379;
  LPM_q_ivl_13359 <= tmp_ivl_13361 & tmp_ivl_13356;
  new_AGEMA_signal_3940 <= tmp_ivl_13363(1);
  n3767 <= tmp_ivl_13363(0);
  tmp_ivl_13363 <= LPM_d0_ivl_13367(0 + 1 downto 0);
  tmp_ivl_13368 <= new_AGEMA_signal_3911 & n3502;
  LPM_q_ivl_13371 <= tmp_ivl_13373 & tmp_ivl_13368;
  tmp_ivl_13375 <= new_AGEMA_signal_3940 & n3767;
  LPM_q_ivl_13378 <= tmp_ivl_13380 & tmp_ivl_13375;
  new_AGEMA_signal_4241 <= tmp_ivl_13382(1);
  n3383 <= tmp_ivl_13382(0);
  tmp_ivl_13382 <= LPM_d0_ivl_13386(0 + 1 downto 0);
  tmp_ivl_13388 <= z1(31);
  tmp_ivl_13389 <= new_AGEMA_signal_3012 & tmp_ivl_13388;
  LPM_q_ivl_13392 <= tmp_ivl_13394 & tmp_ivl_13389;
  tmp_ivl_13397 <= state_in_s1(295);
  tmp_ivl_13399 <= state_in_s0(295);
  tmp_ivl_13400 <= tmp_ivl_13397 & tmp_ivl_13399;
  LPM_q_ivl_13403 <= tmp_ivl_13405 & tmp_ivl_13400;
  new_AGEMA_signal_3379 <= tmp_ivl_13407(1);
  n3382 <= tmp_ivl_13407(0);
  tmp_ivl_13407 <= LPM_d0_ivl_13411(0 + 1 downto 0);
  tmp_ivl_13413 <= z0(31);
  tmp_ivl_13414 <= new_AGEMA_signal_3254 & tmp_ivl_13413;
  LPM_q_ivl_13417 <= tmp_ivl_13419 & tmp_ivl_13414;
  tmp_ivl_13422 <= state_in_s1(39);
  tmp_ivl_13424 <= state_in_s0(39);
  tmp_ivl_13425 <= tmp_ivl_13422 & tmp_ivl_13424;
  LPM_q_ivl_13428 <= tmp_ivl_13430 & tmp_ivl_13425;
  new_AGEMA_signal_3380 <= tmp_ivl_13432(1);
  n3552 <= tmp_ivl_13432(0);
  tmp_ivl_13432 <= LPM_d0_ivl_13436(0 + 1 downto 0);
  tmp_ivl_13438 <= state_in_s1(103);
  tmp_ivl_13440 <= state_in_s0(103);
  tmp_ivl_13441 <= tmp_ivl_13438 & tmp_ivl_13440;
  LPM_q_ivl_13444 <= tmp_ivl_13446 & tmp_ivl_13441;
  tmp_ivl_13448 <= new_AGEMA_signal_3380 & n3552;
  LPM_q_ivl_13451 <= tmp_ivl_13453 & tmp_ivl_13448;
  new_AGEMA_signal_3657 <= tmp_ivl_13455(1);
  n3381 <= tmp_ivl_13455(0);
  tmp_ivl_13455 <= LPM_d0_ivl_13459(0 + 1 downto 0);
  tmp_ivl_13460 <= new_AGEMA_signal_3379 & n3382;
  LPM_q_ivl_13463 <= tmp_ivl_13465 & tmp_ivl_13460;
  tmp_ivl_13467 <= new_AGEMA_signal_3657 & n3381;
  LPM_q_ivl_13470 <= tmp_ivl_13472 & tmp_ivl_13467;
  new_AGEMA_signal_3941 <= tmp_ivl_13474(1);
  n3762 <= tmp_ivl_13474(0);
  tmp_ivl_13474 <= LPM_d0_ivl_13478(0 + 1 downto 0);
  tmp_ivl_13479 <= new_AGEMA_signal_4241 & n3383;
  LPM_q_ivl_13482 <= tmp_ivl_13484 & tmp_ivl_13479;
  tmp_ivl_13486 <= new_AGEMA_signal_3941 & n3762;
  LPM_q_ivl_13489 <= tmp_ivl_13491 & tmp_ivl_13486;
  tmp_ivl_13493 <= tmp_ivl_13497(1);
  tmp_ivl_13495 <= tmp_ivl_13497(0);
  tmp_ivl_13497 <= LPM_d0_ivl_13501(0 + 1 downto 0);
  tmp_ivl_13503 <= z1(26);
  tmp_ivl_13504 <= new_AGEMA_signal_3007 & tmp_ivl_13503;
  LPM_q_ivl_13507 <= tmp_ivl_13509 & tmp_ivl_13504;
  tmp_ivl_13512 <= state_in_s1(290);
  tmp_ivl_13514 <= state_in_s0(290);
  tmp_ivl_13515 <= tmp_ivl_13512 & tmp_ivl_13514;
  LPM_q_ivl_13518 <= tmp_ivl_13520 & tmp_ivl_13515;
  new_AGEMA_signal_3381 <= tmp_ivl_13522(1);
  n3385 <= tmp_ivl_13522(0);
  tmp_ivl_13522 <= LPM_d0_ivl_13526(0 + 1 downto 0);
  tmp_ivl_13528 <= z0(26);
  tmp_ivl_13529 <= new_AGEMA_signal_3258 & tmp_ivl_13528;
  LPM_q_ivl_13532 <= tmp_ivl_13534 & tmp_ivl_13529;
  tmp_ivl_13537 <= state_in_s1(34);
  tmp_ivl_13539 <= state_in_s0(34);
  tmp_ivl_13540 <= tmp_ivl_13537 & tmp_ivl_13539;
  LPM_q_ivl_13543 <= tmp_ivl_13545 & tmp_ivl_13540;
  new_AGEMA_signal_3382 <= tmp_ivl_13547(1);
  n3770 <= tmp_ivl_13547(0);
  tmp_ivl_13547 <= LPM_d0_ivl_13551(0 + 1 downto 0);
  tmp_ivl_13553 <= state_in_s1(98);
  tmp_ivl_13555 <= state_in_s0(98);
  tmp_ivl_13556 <= tmp_ivl_13553 & tmp_ivl_13555;
  LPM_q_ivl_13559 <= tmp_ivl_13561 & tmp_ivl_13556;
  tmp_ivl_13563 <= new_AGEMA_signal_3382 & n3770;
  LPM_q_ivl_13566 <= tmp_ivl_13568 & tmp_ivl_13563;
  new_AGEMA_signal_3658 <= tmp_ivl_13570(1);
  n3384 <= tmp_ivl_13570(0);
  tmp_ivl_13570 <= LPM_d0_ivl_13574(0 + 1 downto 0);
  tmp_ivl_13575 <= new_AGEMA_signal_3381 & n3385;
  LPM_q_ivl_13578 <= tmp_ivl_13580 & tmp_ivl_13575;
  tmp_ivl_13582 <= new_AGEMA_signal_3658 & n3384;
  LPM_q_ivl_13585 <= tmp_ivl_13587 & tmp_ivl_13582;
  new_AGEMA_signal_3942 <= tmp_ivl_13589(1);
  n3898 <= tmp_ivl_13589(0);
  tmp_ivl_13589 <= LPM_d0_ivl_13593(0 + 1 downto 0);
  tmp_ivl_13595 <= z0(48);
  tmp_ivl_13596 <= new_AGEMA_signal_3238 & tmp_ivl_13595;
  LPM_q_ivl_13599 <= tmp_ivl_13601 & tmp_ivl_13596;
  tmp_ivl_13604 <= state_in_s1(8);
  tmp_ivl_13606 <= state_in_s0(8);
  tmp_ivl_13607 <= tmp_ivl_13604 & tmp_ivl_13606;
  LPM_q_ivl_13610 <= tmp_ivl_13612 & tmp_ivl_13607;
  new_AGEMA_signal_3383 <= tmp_ivl_13614(1);
  n3528 <= tmp_ivl_13614(0);
  tmp_ivl_13614 <= LPM_d0_ivl_13618(0 + 1 downto 0);
  tmp_ivl_13620 <= z1(48);
  tmp_ivl_13621 <= new_AGEMA_signal_3029 & tmp_ivl_13620;
  LPM_q_ivl_13624 <= tmp_ivl_13626 & tmp_ivl_13621;
  tmp_ivl_13628 <= new_AGEMA_signal_3383 & n3528;
  LPM_q_ivl_13631 <= tmp_ivl_13633 & tmp_ivl_13628;
  new_AGEMA_signal_3659 <= tmp_ivl_13635(1);
  n3387 <= tmp_ivl_13635(0);
  tmp_ivl_13635 <= LPM_d0_ivl_13639(0 + 1 downto 0);
  tmp_ivl_13640 <= new_AGEMA_signal_3659 & n3387;
  LPM_q_ivl_13643 <= tmp_ivl_13645 & tmp_ivl_13640;
  tmp_ivl_13647 <= new_AGEMA_signal_2671 & n3386;
  LPM_q_ivl_13650 <= tmp_ivl_13652 & tmp_ivl_13647;
  new_AGEMA_signal_3943 <= tmp_ivl_13654(1);
  n3791 <= tmp_ivl_13654(0);
  tmp_ivl_13654 <= LPM_d0_ivl_13658(0 + 1 downto 0);
  tmp_ivl_13659 <= new_AGEMA_signal_3942 & n3898;
  LPM_q_ivl_13662 <= tmp_ivl_13664 & tmp_ivl_13659;
  tmp_ivl_13666 <= new_AGEMA_signal_3943 & n3791;
  LPM_q_ivl_13669 <= tmp_ivl_13671 & tmp_ivl_13666;
  new_AGEMA_signal_4242 <= tmp_ivl_13673(1);
  n3390 <= tmp_ivl_13673(0);
  tmp_ivl_13673 <= LPM_d0_ivl_13677(0 + 1 downto 0);
  tmp_ivl_13679 <= z0(51);
  tmp_ivl_13680 <= new_AGEMA_signal_3234 & tmp_ivl_13679;
  LPM_q_ivl_13683 <= tmp_ivl_13685 & tmp_ivl_13680;
  tmp_ivl_13688 <= state_in_s1(11);
  tmp_ivl_13690 <= state_in_s0(11);
  tmp_ivl_13691 <= tmp_ivl_13688 & tmp_ivl_13690;
  LPM_q_ivl_13694 <= tmp_ivl_13696 & tmp_ivl_13691;
  new_AGEMA_signal_3384 <= tmp_ivl_13698(1);
  n3824 <= tmp_ivl_13698(0);
  tmp_ivl_13698 <= LPM_d0_ivl_13702(0 + 1 downto 0);
  tmp_ivl_13704 <= z1(51);
  tmp_ivl_13705 <= new_AGEMA_signal_3032 & tmp_ivl_13704;
  LPM_q_ivl_13708 <= tmp_ivl_13710 & tmp_ivl_13705;
  tmp_ivl_13712 <= new_AGEMA_signal_3384 & n3824;
  LPM_q_ivl_13715 <= tmp_ivl_13717 & tmp_ivl_13712;
  new_AGEMA_signal_3660 <= tmp_ivl_13719(1);
  n3389 <= tmp_ivl_13719(0);
  tmp_ivl_13719 <= LPM_d0_ivl_13723(0 + 1 downto 0);
  tmp_ivl_13724 <= new_AGEMA_signal_3660 & n3389;
  LPM_q_ivl_13727 <= tmp_ivl_13729 & tmp_ivl_13724;
  tmp_ivl_13731 <= new_AGEMA_signal_2673 & n3388;
  LPM_q_ivl_13734 <= tmp_ivl_13736 & tmp_ivl_13731;
  new_AGEMA_signal_3944 <= tmp_ivl_13738(1);
  n3519 <= tmp_ivl_13738(0);
  tmp_ivl_13738 <= LPM_d0_ivl_13742(0 + 1 downto 0);
  tmp_ivl_13743 <= new_AGEMA_signal_4242 & n3390;
  LPM_q_ivl_13746 <= tmp_ivl_13748 & tmp_ivl_13743;
  tmp_ivl_13750 <= new_AGEMA_signal_3944 & n3519;
  LPM_q_ivl_13753 <= tmp_ivl_13755 & tmp_ivl_13750;
  tmp_ivl_13757 <= tmp_ivl_13761(1);
  tmp_ivl_13759 <= tmp_ivl_13761(0);
  tmp_ivl_13761 <= LPM_d0_ivl_13765(0 + 1 downto 0);
  tmp_ivl_13766 <= new_AGEMA_signal_3596 & n3391;
  LPM_q_ivl_13769 <= tmp_ivl_13771 & tmp_ivl_13766;
  tmp_ivl_13773 <= new_AGEMA_signal_3618 & n3629;
  LPM_q_ivl_13776 <= tmp_ivl_13778 & tmp_ivl_13773;
  new_AGEMA_signal_3945 <= tmp_ivl_13780(1);
  n3392 <= tmp_ivl_13780(0);
  tmp_ivl_13780 <= LPM_d0_ivl_13784(0 + 1 downto 0);
  tmp_ivl_13786 <= state_in_s1(196);
  tmp_ivl_13788 <= state_in_s0(196);
  tmp_ivl_13789 <= tmp_ivl_13786 & tmp_ivl_13788;
  LPM_q_ivl_13792 <= tmp_ivl_13794 & tmp_ivl_13789;
  tmp_ivl_13797 <= z4(60);
  tmp_ivl_13798 <= new_AGEMA_signal_3167 & tmp_ivl_13797;
  LPM_q_ivl_13801 <= tmp_ivl_13803 & tmp_ivl_13798;
  new_AGEMA_signal_3385 <= tmp_ivl_13805(1);
  n3485 <= tmp_ivl_13805(0);
  tmp_ivl_13805 <= LPM_d0_ivl_13809(0 + 1 downto 0);
  tmp_ivl_13811 <= state_in_s1(260);
  tmp_ivl_13813 <= state_in_s0(260);
  tmp_ivl_13814 <= tmp_ivl_13811 & tmp_ivl_13813;
  LPM_q_ivl_13817 <= tmp_ivl_13819 & tmp_ivl_13814;
  tmp_ivl_13821 <= new_AGEMA_signal_3385 & n3485;
  LPM_q_ivl_13824 <= tmp_ivl_13826 & tmp_ivl_13821;
  new_AGEMA_signal_3661 <= tmp_ivl_13828(1);
  n3624 <= tmp_ivl_13828(0);
  tmp_ivl_13828 <= LPM_d0_ivl_13832(0 + 1 downto 0);
  tmp_ivl_13833 <= new_AGEMA_signal_3945 & n3392;
  LPM_q_ivl_13836 <= tmp_ivl_13838 & tmp_ivl_13833;
  tmp_ivl_13840 <= new_AGEMA_signal_3661 & n3624;
  LPM_q_ivl_13843 <= tmp_ivl_13845 & tmp_ivl_13840;
  tmp_ivl_13847 <= tmp_ivl_13851(1);
  tmp_ivl_13849 <= tmp_ivl_13851(0);
  tmp_ivl_13851 <= LPM_d0_ivl_13855(0 + 1 downto 0);
  tmp_ivl_13856 <= new_AGEMA_signal_3600 & n3660;
  LPM_q_ivl_13859 <= tmp_ivl_13861 & tmp_ivl_13856;
  tmp_ivl_13863 <= new_AGEMA_signal_3654 & n3656;
  LPM_q_ivl_13866 <= tmp_ivl_13868 & tmp_ivl_13863;
  new_AGEMA_signal_3946 <= tmp_ivl_13870(1);
  n3393 <= tmp_ivl_13870(0);
  tmp_ivl_13870 <= LPM_d0_ivl_13874(0 + 1 downto 0);
  tmp_ivl_13875 <= new_AGEMA_signal_3946 & n3393;
  LPM_q_ivl_13878 <= tmp_ivl_13880 & tmp_ivl_13875;
  tmp_ivl_13882 <= new_AGEMA_signal_3661 & n3624;
  LPM_q_ivl_13885 <= tmp_ivl_13887 & tmp_ivl_13882;
  tmp_ivl_13889 <= tmp_ivl_13893(1);
  tmp_ivl_13891 <= tmp_ivl_13893(0);
  tmp_ivl_13893 <= LPM_d0_ivl_13897(0 + 1 downto 0);
  tmp_ivl_13898 <= new_AGEMA_signal_3336 & n3395;
  LPM_q_ivl_13901 <= tmp_ivl_13903 & tmp_ivl_13898;
  tmp_ivl_13905 <= new_AGEMA_signal_3331 & n3394;
  LPM_q_ivl_13908 <= tmp_ivl_13910 & tmp_ivl_13905;
  new_AGEMA_signal_3662 <= tmp_ivl_13912(1);
  n3846 <= tmp_ivl_13912(0);
  tmp_ivl_13912 <= LPM_d0_ivl_13916(0 + 1 downto 0);
  tmp_ivl_13917 <= new_AGEMA_signal_3645 & n3637;
  LPM_q_ivl_13920 <= tmp_ivl_13922 & tmp_ivl_13917;
  tmp_ivl_13924 <= new_AGEMA_signal_3662 & n3846;
  LPM_q_ivl_13927 <= tmp_ivl_13929 & tmp_ivl_13924;
  new_AGEMA_signal_3947 <= tmp_ivl_13931(1);
  n3397 <= tmp_ivl_13931(0);
  tmp_ivl_13931 <= LPM_d0_ivl_13935(0 + 1 downto 0);
  tmp_ivl_13937 <= z0(10);
  tmp_ivl_13938 <= new_AGEMA_signal_3230 & tmp_ivl_13937;
  LPM_q_ivl_13941 <= tmp_ivl_13943 & tmp_ivl_13938;
  tmp_ivl_13946 <= state_in_s1(50);
  tmp_ivl_13948 <= state_in_s0(50);
  tmp_ivl_13949 <= tmp_ivl_13946 & tmp_ivl_13948;
  LPM_q_ivl_13952 <= tmp_ivl_13954 & tmp_ivl_13949;
  new_AGEMA_signal_3386 <= tmp_ivl_13956(1);
  n3398 <= tmp_ivl_13956(0);
  tmp_ivl_13956 <= LPM_d0_ivl_13960(0 + 1 downto 0);
  tmp_ivl_13961 <= new_AGEMA_signal_3386 & n3398;
  LPM_q_ivl_13964 <= tmp_ivl_13966 & tmp_ivl_13961;
  tmp_ivl_13968 <= new_AGEMA_signal_3304 & n3396;
  LPM_q_ivl_13971 <= tmp_ivl_13973 & tmp_ivl_13968;
  new_AGEMA_signal_3663 <= tmp_ivl_13975(1);
  n3843 <= tmp_ivl_13975(0);
  tmp_ivl_13975 <= LPM_d0_ivl_13979(0 + 1 downto 0);
  tmp_ivl_13980 <= new_AGEMA_signal_3947 & n3397;
  LPM_q_ivl_13983 <= tmp_ivl_13985 & tmp_ivl_13980;
  tmp_ivl_13987 <= new_AGEMA_signal_3663 & n3843;
  LPM_q_ivl_13990 <= tmp_ivl_13992 & tmp_ivl_13987;
  tmp_ivl_13994 <= tmp_ivl_13998(1);
  tmp_ivl_13996 <= tmp_ivl_13998(0);
  tmp_ivl_13998 <= LPM_d0_ivl_14002(0 + 1 downto 0);
  tmp_ivl_14004 <= z1(10);
  tmp_ivl_14005 <= new_AGEMA_signal_2991 & tmp_ivl_14004;
  LPM_q_ivl_14008 <= tmp_ivl_14010 & tmp_ivl_14005;
  tmp_ivl_14013 <= state_in_s1(306);
  tmp_ivl_14015 <= state_in_s0(306);
  tmp_ivl_14016 <= tmp_ivl_14013 & tmp_ivl_14015;
  LPM_q_ivl_14019 <= tmp_ivl_14021 & tmp_ivl_14016;
  new_AGEMA_signal_3387 <= tmp_ivl_14023(1);
  n3400 <= tmp_ivl_14023(0);
  tmp_ivl_14023 <= LPM_d0_ivl_14027(0 + 1 downto 0);
  tmp_ivl_14029 <= state_in_s1(114);
  tmp_ivl_14031 <= state_in_s0(114);
  tmp_ivl_14032 <= tmp_ivl_14029 & tmp_ivl_14031;
  LPM_q_ivl_14035 <= tmp_ivl_14037 & tmp_ivl_14032;
  tmp_ivl_14039 <= new_AGEMA_signal_3386 & n3398;
  LPM_q_ivl_14042 <= tmp_ivl_14044 & tmp_ivl_14039;
  new_AGEMA_signal_3664 <= tmp_ivl_14046(1);
  n3399 <= tmp_ivl_14046(0);
  tmp_ivl_14046 <= LPM_d0_ivl_14050(0 + 1 downto 0);
  tmp_ivl_14051 <= new_AGEMA_signal_3387 & n3400;
  LPM_q_ivl_14054 <= tmp_ivl_14056 & tmp_ivl_14051;
  tmp_ivl_14058 <= new_AGEMA_signal_3664 & n3399;
  LPM_q_ivl_14061 <= tmp_ivl_14063 & tmp_ivl_14058;
  new_AGEMA_signal_3948 <= tmp_ivl_14065(1);
  n3884 <= tmp_ivl_14065(0);
  tmp_ivl_14065 <= LPM_d0_ivl_14069(0 + 1 downto 0);
  tmp_ivl_14070 <= new_AGEMA_signal_3918 & n3412;
  LPM_q_ivl_14073 <= tmp_ivl_14075 & tmp_ivl_14070;
  tmp_ivl_14077 <= new_AGEMA_signal_3948 & n3884;
  LPM_q_ivl_14080 <= tmp_ivl_14082 & tmp_ivl_14077;
  new_AGEMA_signal_4246 <= tmp_ivl_14084(1);
  n3403 <= tmp_ivl_14084(0);
  tmp_ivl_14084 <= LPM_d0_ivl_14088(0 + 1 downto 0);
  tmp_ivl_14090 <= z1(32);
  tmp_ivl_14091 <= new_AGEMA_signal_3013 & tmp_ivl_14090;
  LPM_q_ivl_14094 <= tmp_ivl_14096 & tmp_ivl_14091;
  tmp_ivl_14099 <= state_in_s1(280);
  tmp_ivl_14101 <= state_in_s0(280);
  tmp_ivl_14102 <= tmp_ivl_14099 & tmp_ivl_14101;
  LPM_q_ivl_14105 <= tmp_ivl_14107 & tmp_ivl_14102;
  new_AGEMA_signal_3388 <= tmp_ivl_14109(1);
  n3402 <= tmp_ivl_14109(0);
  tmp_ivl_14109 <= LPM_d0_ivl_14113(0 + 1 downto 0);
  tmp_ivl_14115 <= z0(32);
  tmp_ivl_14116 <= new_AGEMA_signal_3268 & tmp_ivl_14115;
  LPM_q_ivl_14119 <= tmp_ivl_14121 & tmp_ivl_14116;
  tmp_ivl_14124 <= state_in_s1(24);
  tmp_ivl_14126 <= state_in_s0(24);
  tmp_ivl_14127 <= tmp_ivl_14124 & tmp_ivl_14126;
  LPM_q_ivl_14130 <= tmp_ivl_14132 & tmp_ivl_14127;
  new_AGEMA_signal_3389 <= tmp_ivl_14134(1);
  n3604 <= tmp_ivl_14134(0);
  tmp_ivl_14134 <= LPM_d0_ivl_14138(0 + 1 downto 0);
  tmp_ivl_14140 <= state_in_s1(88);
  tmp_ivl_14142 <= state_in_s0(88);
  tmp_ivl_14143 <= tmp_ivl_14140 & tmp_ivl_14142;
  LPM_q_ivl_14146 <= tmp_ivl_14148 & tmp_ivl_14143;
  tmp_ivl_14150 <= new_AGEMA_signal_3389 & n3604;
  LPM_q_ivl_14153 <= tmp_ivl_14155 & tmp_ivl_14150;
  new_AGEMA_signal_3665 <= tmp_ivl_14157(1);
  n3401 <= tmp_ivl_14157(0);
  tmp_ivl_14157 <= LPM_d0_ivl_14161(0 + 1 downto 0);
  tmp_ivl_14162 <= new_AGEMA_signal_3388 & n3402;
  LPM_q_ivl_14165 <= tmp_ivl_14167 & tmp_ivl_14162;
  tmp_ivl_14169 <= new_AGEMA_signal_3665 & n3401;
  LPM_q_ivl_14172 <= tmp_ivl_14174 & tmp_ivl_14169;
  new_AGEMA_signal_3949 <= tmp_ivl_14176(1);
  n3878 <= tmp_ivl_14176(0);
  tmp_ivl_14176 <= LPM_d0_ivl_14180(0 + 1 downto 0);
  tmp_ivl_14181 <= new_AGEMA_signal_4246 & n3403;
  LPM_q_ivl_14184 <= tmp_ivl_14186 & tmp_ivl_14181;
  tmp_ivl_14188 <= new_AGEMA_signal_3949 & n3878;
  LPM_q_ivl_14191 <= tmp_ivl_14193 & tmp_ivl_14188;
  tmp_ivl_14195 <= tmp_ivl_14199(1);
  tmp_ivl_14197 <= tmp_ivl_14199(0);
  tmp_ivl_14199 <= LPM_d0_ivl_14203(0 + 1 downto 0);
  tmp_ivl_14205 <= z0(13);
  tmp_ivl_14206 <= new_AGEMA_signal_3231 & tmp_ivl_14205;
  LPM_q_ivl_14209 <= tmp_ivl_14211 & tmp_ivl_14206;
  tmp_ivl_14214 <= state_in_s1(53);
  tmp_ivl_14216 <= state_in_s0(53);
  tmp_ivl_14217 <= tmp_ivl_14214 & tmp_ivl_14216;
  LPM_q_ivl_14220 <= tmp_ivl_14222 & tmp_ivl_14217;
  new_AGEMA_signal_3390 <= tmp_ivl_14224(1);
  n3413 <= tmp_ivl_14224(0);
  tmp_ivl_14224 <= LPM_d0_ivl_14228(0 + 1 downto 0);
  tmp_ivl_14229 <= new_AGEMA_signal_3390 & n3413;
  LPM_q_ivl_14232 <= tmp_ivl_14234 & tmp_ivl_14229;
  tmp_ivl_14236 <= new_AGEMA_signal_3317 & n3404;
  LPM_q_ivl_14239 <= tmp_ivl_14241 & tmp_ivl_14236;
  new_AGEMA_signal_3666 <= tmp_ivl_14243(1);
  n3887 <= tmp_ivl_14243(0);
  tmp_ivl_14243 <= LPM_d0_ivl_14247(0 + 1 downto 0);
  tmp_ivl_14249 <= z0(22);
  tmp_ivl_14250 <= new_AGEMA_signal_3243 & tmp_ivl_14249;
  LPM_q_ivl_14253 <= tmp_ivl_14255 & tmp_ivl_14250;
  tmp_ivl_14258 <= state_in_s1(46);
  tmp_ivl_14260 <= state_in_s0(46);
  tmp_ivl_14261 <= tmp_ivl_14258 & tmp_ivl_14260;
  LPM_q_ivl_14264 <= tmp_ivl_14266 & tmp_ivl_14261;
  new_AGEMA_signal_3391 <= tmp_ivl_14268(1);
  n3546 <= tmp_ivl_14268(0);
  tmp_ivl_14268 <= LPM_d0_ivl_14272(0 + 1 downto 0);
  tmp_ivl_14273 <= new_AGEMA_signal_3391 & n3546;
  LPM_q_ivl_14276 <= tmp_ivl_14278 & tmp_ivl_14273;
  tmp_ivl_14280 <= new_AGEMA_signal_3295 & n3405;
  LPM_q_ivl_14283 <= tmp_ivl_14285 & tmp_ivl_14280;
  new_AGEMA_signal_3667 <= tmp_ivl_14287(1);
  n3806 <= tmp_ivl_14287(0);
  tmp_ivl_14287 <= LPM_d0_ivl_14291(0 + 1 downto 0);
  tmp_ivl_14292 <= new_AGEMA_signal_3666 & n3887;
  LPM_q_ivl_14295 <= tmp_ivl_14297 & tmp_ivl_14292;
  tmp_ivl_14299 <= new_AGEMA_signal_3667 & n3806;
  LPM_q_ivl_14302 <= tmp_ivl_14304 & tmp_ivl_14299;
  new_AGEMA_signal_3950 <= tmp_ivl_14306(1);
  n3408 <= tmp_ivl_14306(0);
  tmp_ivl_14306 <= LPM_d0_ivl_14310(0 + 1 downto 0);
  tmp_ivl_14311 <= new_AGEMA_signal_3332 & n3407;
  LPM_q_ivl_14314 <= tmp_ivl_14316 & tmp_ivl_14311;
  tmp_ivl_14318 <= new_AGEMA_signal_3362 & n3406;
  LPM_q_ivl_14321 <= tmp_ivl_14323 & tmp_ivl_14318;
  new_AGEMA_signal_3668 <= tmp_ivl_14325(1);
  n3803 <= tmp_ivl_14325(0);
  tmp_ivl_14325 <= LPM_d0_ivl_14329(0 + 1 downto 0);
  tmp_ivl_14330 <= new_AGEMA_signal_3950 & n3408;
  LPM_q_ivl_14333 <= tmp_ivl_14335 & tmp_ivl_14330;
  tmp_ivl_14337 <= new_AGEMA_signal_3668 & n3803;
  LPM_q_ivl_14340 <= tmp_ivl_14342 & tmp_ivl_14337;
  tmp_ivl_14344 <= tmp_ivl_14348(1);
  tmp_ivl_14346 <= tmp_ivl_14348(0);
  tmp_ivl_14348 <= LPM_d0_ivl_14352(0 + 1 downto 0);
  tmp_ivl_14354 <= z1(38);
  tmp_ivl_14355 <= new_AGEMA_signal_3019 & tmp_ivl_14354;
  LPM_q_ivl_14358 <= tmp_ivl_14360 & tmp_ivl_14355;
  tmp_ivl_14363 <= state_in_s1(286);
  tmp_ivl_14365 <= state_in_s0(286);
  tmp_ivl_14366 <= tmp_ivl_14363 & tmp_ivl_14365;
  LPM_q_ivl_14369 <= tmp_ivl_14371 & tmp_ivl_14366;
  new_AGEMA_signal_3392 <= tmp_ivl_14373(1);
  n3411 <= tmp_ivl_14373(0);
  tmp_ivl_14373 <= LPM_d0_ivl_14377(0 + 1 downto 0);
  tmp_ivl_14379 <= state_in_s1(94);
  tmp_ivl_14381 <= state_in_s0(94);
  tmp_ivl_14382 <= tmp_ivl_14379 & tmp_ivl_14381;
  LPM_q_ivl_14385 <= tmp_ivl_14387 & tmp_ivl_14382;
  tmp_ivl_14389 <= new_AGEMA_signal_3363 & n3409;
  LPM_q_ivl_14392 <= tmp_ivl_14394 & tmp_ivl_14389;
  new_AGEMA_signal_3669 <= tmp_ivl_14396(1);
  n3410 <= tmp_ivl_14396(0);
  tmp_ivl_14396 <= LPM_d0_ivl_14400(0 + 1 downto 0);
  tmp_ivl_14401 <= new_AGEMA_signal_3392 & n3411;
  LPM_q_ivl_14404 <= tmp_ivl_14406 & tmp_ivl_14401;
  tmp_ivl_14408 <= new_AGEMA_signal_3669 & n3410;
  LPM_q_ivl_14411 <= tmp_ivl_14413 & tmp_ivl_14408;
  new_AGEMA_signal_3951 <= tmp_ivl_14415(1);
  n3607 <= tmp_ivl_14415(0);
  tmp_ivl_14415 <= LPM_d0_ivl_14419(0 + 1 downto 0);
  tmp_ivl_14420 <= new_AGEMA_signal_3918 & n3412;
  LPM_q_ivl_14423 <= tmp_ivl_14425 & tmp_ivl_14420;
  tmp_ivl_14427 <= new_AGEMA_signal_3951 & n3607;
  LPM_q_ivl_14430 <= tmp_ivl_14432 & tmp_ivl_14427;
  new_AGEMA_signal_4248 <= tmp_ivl_14434(1);
  n3416 <= tmp_ivl_14434(0);
  tmp_ivl_14434 <= LPM_d0_ivl_14438(0 + 1 downto 0);
  tmp_ivl_14440 <= z1(13);
  tmp_ivl_14441 <= new_AGEMA_signal_2994 & tmp_ivl_14440;
  LPM_q_ivl_14444 <= tmp_ivl_14446 & tmp_ivl_14441;
  tmp_ivl_14449 <= state_in_s1(309);
  tmp_ivl_14451 <= state_in_s0(309);
  tmp_ivl_14452 <= tmp_ivl_14449 & tmp_ivl_14451;
  LPM_q_ivl_14455 <= tmp_ivl_14457 & tmp_ivl_14452;
  new_AGEMA_signal_3393 <= tmp_ivl_14459(1);
  n3415 <= tmp_ivl_14459(0);
  tmp_ivl_14459 <= LPM_d0_ivl_14463(0 + 1 downto 0);
  tmp_ivl_14465 <= state_in_s1(117);
  tmp_ivl_14467 <= state_in_s0(117);
  tmp_ivl_14468 <= tmp_ivl_14465 & tmp_ivl_14467;
  LPM_q_ivl_14471 <= tmp_ivl_14473 & tmp_ivl_14468;
  tmp_ivl_14475 <= new_AGEMA_signal_3390 & n3413;
  LPM_q_ivl_14478 <= tmp_ivl_14480 & tmp_ivl_14475;
  new_AGEMA_signal_3670 <= tmp_ivl_14482(1);
  n3414 <= tmp_ivl_14482(0);
  tmp_ivl_14482 <= LPM_d0_ivl_14486(0 + 1 downto 0);
  tmp_ivl_14487 <= new_AGEMA_signal_3393 & n3415;
  LPM_q_ivl_14490 <= tmp_ivl_14492 & tmp_ivl_14487;
  tmp_ivl_14494 <= new_AGEMA_signal_3670 & n3414;
  LPM_q_ivl_14497 <= tmp_ivl_14499 & tmp_ivl_14494;
  new_AGEMA_signal_3952 <= tmp_ivl_14501(1);
  n3435 <= tmp_ivl_14501(0);
  tmp_ivl_14501 <= LPM_d0_ivl_14505(0 + 1 downto 0);
  tmp_ivl_14506 <= new_AGEMA_signal_4248 & n3416;
  LPM_q_ivl_14509 <= tmp_ivl_14511 & tmp_ivl_14506;
  tmp_ivl_14513 <= new_AGEMA_signal_3952 & n3435;
  LPM_q_ivl_14516 <= tmp_ivl_14518 & tmp_ivl_14513;
  tmp_ivl_14520 <= tmp_ivl_14524(1);
  tmp_ivl_14522 <= tmp_ivl_14524(0);
  tmp_ivl_14524 <= LPM_d0_ivl_14528(0 + 1 downto 0);
  tmp_ivl_14529 <= new_AGEMA_signal_3909 & n3433;
  LPM_q_ivl_14532 <= tmp_ivl_14534 & tmp_ivl_14529;
  tmp_ivl_14536 <= new_AGEMA_signal_3922 & n3608;
  LPM_q_ivl_14539 <= tmp_ivl_14541 & tmp_ivl_14536;
  new_AGEMA_signal_4249 <= tmp_ivl_14543(1);
  n3417 <= tmp_ivl_14543(0);
  tmp_ivl_14543 <= LPM_d0_ivl_14547(0 + 1 downto 0);
  tmp_ivl_14548 <= new_AGEMA_signal_4249 & n3417;
  LPM_q_ivl_14551 <= tmp_ivl_14553 & tmp_ivl_14548;
  tmp_ivl_14555 <= new_AGEMA_signal_3952 & n3435;
  LPM_q_ivl_14558 <= tmp_ivl_14560 & tmp_ivl_14555;
  tmp_ivl_14562 <= tmp_ivl_14566(1);
  tmp_ivl_14564 <= tmp_ivl_14566(0);
  tmp_ivl_14566 <= LPM_d0_ivl_14570(0 + 1 downto 0);
  tmp_ivl_14572 <= z0(27);
  tmp_ivl_14573 <= new_AGEMA_signal_3257 & tmp_ivl_14572;
  LPM_q_ivl_14576 <= tmp_ivl_14578 & tmp_ivl_14573;
  tmp_ivl_14581 <= state_in_s1(35);
  tmp_ivl_14583 <= state_in_s0(35);
  tmp_ivl_14584 <= tmp_ivl_14581 & tmp_ivl_14583;
  LPM_q_ivl_14587 <= tmp_ivl_14589 & tmp_ivl_14584;
  new_AGEMA_signal_3394 <= tmp_ivl_14591(1);
  n3427 <= tmp_ivl_14591(0);
  tmp_ivl_14591 <= LPM_d0_ivl_14595(0 + 1 downto 0);
  tmp_ivl_14597 <= state_in_s1(227);
  tmp_ivl_14599 <= state_in_s0(227);
  tmp_ivl_14600 <= tmp_ivl_14597 & tmp_ivl_14599;
  LPM_q_ivl_14603 <= tmp_ivl_14605 & tmp_ivl_14600;
  tmp_ivl_14608 <= z4(27);
  tmp_ivl_14609 <= new_AGEMA_signal_3130 & tmp_ivl_14608;
  LPM_q_ivl_14612 <= tmp_ivl_14614 & tmp_ivl_14609;
  new_AGEMA_signal_3395 <= tmp_ivl_14616(1);
  n3423 <= tmp_ivl_14616(0);
  tmp_ivl_14616 <= LPM_d0_ivl_14620(0 + 1 downto 0);
  tmp_ivl_14621 <= new_AGEMA_signal_3394 & n3427;
  LPM_q_ivl_14624 <= tmp_ivl_14626 & tmp_ivl_14621;
  tmp_ivl_14628 <= new_AGEMA_signal_3395 & n3423;
  LPM_q_ivl_14631 <= tmp_ivl_14633 & tmp_ivl_14628;
  new_AGEMA_signal_3671 <= tmp_ivl_14635(1);
  n3856 <= tmp_ivl_14635(0);
  tmp_ivl_14635 <= LPM_d0_ivl_14639(0 + 1 downto 0);
  tmp_ivl_14641 <= z0(36);
  tmp_ivl_14642 <= new_AGEMA_signal_3262 & tmp_ivl_14641;
  LPM_q_ivl_14645 <= tmp_ivl_14647 & tmp_ivl_14642;
  tmp_ivl_14650 <= state_in_s1(28);
  tmp_ivl_14652 <= state_in_s0(28);
  tmp_ivl_14653 <= tmp_ivl_14650 & tmp_ivl_14652;
  LPM_q_ivl_14656 <= tmp_ivl_14658 & tmp_ivl_14653;
  new_AGEMA_signal_3396 <= tmp_ivl_14660(1);
  n3444 <= tmp_ivl_14660(0);
  tmp_ivl_14660 <= LPM_d0_ivl_14664(0 + 1 downto 0);
  tmp_ivl_14665 <= new_AGEMA_signal_3396 & n3444;
  LPM_q_ivl_14668 <= tmp_ivl_14670 & tmp_ivl_14665;
  tmp_ivl_14672 <= new_AGEMA_signal_3327 & n3418;
  LPM_q_ivl_14675 <= tmp_ivl_14677 & tmp_ivl_14672;
  new_AGEMA_signal_3672 <= tmp_ivl_14679(1);
  n3787 <= tmp_ivl_14679(0);
  tmp_ivl_14679 <= LPM_d0_ivl_14683(0 + 1 downto 0);
  tmp_ivl_14684 <= new_AGEMA_signal_3671 & n3856;
  LPM_q_ivl_14687 <= tmp_ivl_14689 & tmp_ivl_14684;
  tmp_ivl_14691 <= new_AGEMA_signal_3672 & n3787;
  LPM_q_ivl_14694 <= tmp_ivl_14696 & tmp_ivl_14691;
  new_AGEMA_signal_3953 <= tmp_ivl_14698(1);
  n3421 <= tmp_ivl_14698(0);
  tmp_ivl_14698 <= LPM_d0_ivl_14702(0 + 1 downto 0);
  tmp_ivl_14703 <= new_AGEMA_signal_3369 & n3420;
  LPM_q_ivl_14706 <= tmp_ivl_14708 & tmp_ivl_14703;
  tmp_ivl_14710 <= new_AGEMA_signal_3298 & n3419;
  LPM_q_ivl_14713 <= tmp_ivl_14715 & tmp_ivl_14710;
  new_AGEMA_signal_3673 <= tmp_ivl_14717(1);
  n3774 <= tmp_ivl_14717(0);
  tmp_ivl_14717 <= LPM_d0_ivl_14721(0 + 1 downto 0);
  tmp_ivl_14722 <= new_AGEMA_signal_3953 & n3421;
  LPM_q_ivl_14725 <= tmp_ivl_14727 & tmp_ivl_14722;
  tmp_ivl_14729 <= new_AGEMA_signal_3673 & n3774;
  LPM_q_ivl_14732 <= tmp_ivl_14734 & tmp_ivl_14729;
  tmp_ivl_14736 <= tmp_ivl_14740(1);
  tmp_ivl_14738 <= tmp_ivl_14740(0);
  tmp_ivl_14740 <= LPM_d0_ivl_14744(0 + 1 downto 0);
  tmp_ivl_14745 <= new_AGEMA_signal_3599 & n3454;
  LPM_q_ivl_14748 <= tmp_ivl_14750 & tmp_ivl_14745;
  tmp_ivl_14752 <= new_AGEMA_signal_3615 & n3422;
  LPM_q_ivl_14755 <= tmp_ivl_14757 & tmp_ivl_14752;
  new_AGEMA_signal_3954 <= tmp_ivl_14759(1);
  n3424 <= tmp_ivl_14759(0);
  tmp_ivl_14759 <= LPM_d0_ivl_14763(0 + 1 downto 0);
  tmp_ivl_14765 <= state_in_s1(291);
  tmp_ivl_14767 <= state_in_s0(291);
  tmp_ivl_14768 <= tmp_ivl_14765 & tmp_ivl_14767;
  LPM_q_ivl_14771 <= tmp_ivl_14773 & tmp_ivl_14768;
  tmp_ivl_14775 <= new_AGEMA_signal_3395 & n3423;
  LPM_q_ivl_14778 <= tmp_ivl_14780 & tmp_ivl_14775;
  new_AGEMA_signal_3674 <= tmp_ivl_14782(1);
  n3725 <= tmp_ivl_14782(0);
  tmp_ivl_14782 <= LPM_d0_ivl_14786(0 + 1 downto 0);
  tmp_ivl_14787 <= new_AGEMA_signal_3954 & n3424;
  LPM_q_ivl_14790 <= tmp_ivl_14792 & tmp_ivl_14787;
  tmp_ivl_14794 <= new_AGEMA_signal_3674 & n3725;
  LPM_q_ivl_14797 <= tmp_ivl_14799 & tmp_ivl_14794;
  tmp_ivl_14801 <= tmp_ivl_14805(1);
  tmp_ivl_14803 <= tmp_ivl_14805(0);
  tmp_ivl_14805 <= LPM_d0_ivl_14809(0 + 1 downto 0);
  tmp_ivl_14811 <= z1(49);
  tmp_ivl_14812 <= new_AGEMA_signal_3030 & tmp_ivl_14811;
  LPM_q_ivl_14815 <= tmp_ivl_14817 & tmp_ivl_14812;
  tmp_ivl_14820 <= state_in_s1(265);
  tmp_ivl_14822 <= state_in_s0(265);
  tmp_ivl_14823 <= tmp_ivl_14820 & tmp_ivl_14822;
  LPM_q_ivl_14826 <= tmp_ivl_14828 & tmp_ivl_14823;
  new_AGEMA_signal_3397 <= tmp_ivl_14830(1);
  n3426 <= tmp_ivl_14830(0);
  tmp_ivl_14830 <= LPM_d0_ivl_14834(0 + 1 downto 0);
  tmp_ivl_14836 <= z0(49);
  tmp_ivl_14837 <= new_AGEMA_signal_3237 & tmp_ivl_14836;
  LPM_q_ivl_14840 <= tmp_ivl_14842 & tmp_ivl_14837;
  tmp_ivl_14845 <= state_in_s1(9);
  tmp_ivl_14847 <= state_in_s0(9);
  tmp_ivl_14848 <= tmp_ivl_14845 & tmp_ivl_14847;
  LPM_q_ivl_14851 <= tmp_ivl_14853 & tmp_ivl_14848;
  new_AGEMA_signal_3398 <= tmp_ivl_14855(1);
  n3653 <= tmp_ivl_14855(0);
  tmp_ivl_14855 <= LPM_d0_ivl_14859(0 + 1 downto 0);
  tmp_ivl_14861 <= state_in_s1(73);
  tmp_ivl_14863 <= state_in_s0(73);
  tmp_ivl_14864 <= tmp_ivl_14861 & tmp_ivl_14863;
  LPM_q_ivl_14867 <= tmp_ivl_14869 & tmp_ivl_14864;
  tmp_ivl_14871 <= new_AGEMA_signal_3398 & n3653;
  LPM_q_ivl_14874 <= tmp_ivl_14876 & tmp_ivl_14871;
  new_AGEMA_signal_3675 <= tmp_ivl_14878(1);
  n3425 <= tmp_ivl_14878(0);
  tmp_ivl_14878 <= LPM_d0_ivl_14882(0 + 1 downto 0);
  tmp_ivl_14883 <= new_AGEMA_signal_3397 & n3426;
  LPM_q_ivl_14886 <= tmp_ivl_14888 & tmp_ivl_14883;
  tmp_ivl_14890 <= new_AGEMA_signal_3675 & n3425;
  LPM_q_ivl_14893 <= tmp_ivl_14895 & tmp_ivl_14890;
  new_AGEMA_signal_3955 <= tmp_ivl_14897(1);
  n3883 <= tmp_ivl_14897(0);
  tmp_ivl_14897 <= LPM_d0_ivl_14901(0 + 1 downto 0);
  tmp_ivl_14903 <= z1(27);
  tmp_ivl_14904 <= new_AGEMA_signal_3008 & tmp_ivl_14903;
  LPM_q_ivl_14907 <= tmp_ivl_14909 & tmp_ivl_14904;
  tmp_ivl_14912 <= state_in_s1(291);
  tmp_ivl_14914 <= state_in_s0(291);
  tmp_ivl_14915 <= tmp_ivl_14912 & tmp_ivl_14914;
  LPM_q_ivl_14918 <= tmp_ivl_14920 & tmp_ivl_14915;
  new_AGEMA_signal_3399 <= tmp_ivl_14922(1);
  n3429 <= tmp_ivl_14922(0);
  tmp_ivl_14922 <= LPM_d0_ivl_14926(0 + 1 downto 0);
  tmp_ivl_14928 <= state_in_s1(99);
  tmp_ivl_14930 <= state_in_s0(99);
  tmp_ivl_14931 <= tmp_ivl_14928 & tmp_ivl_14930;
  LPM_q_ivl_14934 <= tmp_ivl_14936 & tmp_ivl_14931;
  tmp_ivl_14938 <= new_AGEMA_signal_3394 & n3427;
  LPM_q_ivl_14941 <= tmp_ivl_14943 & tmp_ivl_14938;
  new_AGEMA_signal_3676 <= tmp_ivl_14945(1);
  n3428 <= tmp_ivl_14945(0);
  tmp_ivl_14945 <= LPM_d0_ivl_14949(0 + 1 downto 0);
  tmp_ivl_14950 <= new_AGEMA_signal_3399 & n3429;
  LPM_q_ivl_14953 <= tmp_ivl_14955 & tmp_ivl_14950;
  tmp_ivl_14957 <= new_AGEMA_signal_3676 & n3428;
  LPM_q_ivl_14960 <= tmp_ivl_14962 & tmp_ivl_14957;
  new_AGEMA_signal_3956 <= tmp_ivl_14964(1);
  n3744 <= tmp_ivl_14964(0);
  tmp_ivl_14964 <= LPM_d0_ivl_14968(0 + 1 downto 0);
  tmp_ivl_14969 <= new_AGEMA_signal_3955 & n3883;
  LPM_q_ivl_14972 <= tmp_ivl_14974 & tmp_ivl_14969;
  tmp_ivl_14976 <= new_AGEMA_signal_3956 & n3744;
  LPM_q_ivl_14979 <= tmp_ivl_14981 & tmp_ivl_14976;
  new_AGEMA_signal_4252 <= tmp_ivl_14983(1);
  n3432 <= tmp_ivl_14983(0);
  tmp_ivl_14983 <= LPM_d0_ivl_14987(0 + 1 downto 0);
  tmp_ivl_14989 <= z0(52);
  tmp_ivl_14990 <= new_AGEMA_signal_3232 & tmp_ivl_14989;
  LPM_q_ivl_14993 <= tmp_ivl_14995 & tmp_ivl_14990;
  tmp_ivl_14998 <= state_in_s1(12);
  tmp_ivl_15000 <= state_in_s0(12);
  tmp_ivl_15001 <= tmp_ivl_14998 & tmp_ivl_15000;
  LPM_q_ivl_15004 <= tmp_ivl_15006 & tmp_ivl_15001;
  new_AGEMA_signal_3400 <= tmp_ivl_15008(1);
  n3912 <= tmp_ivl_15008(0);
  tmp_ivl_15008 <= LPM_d0_ivl_15012(0 + 1 downto 0);
  tmp_ivl_15014 <= z1(52);
  tmp_ivl_15015 <= new_AGEMA_signal_3033 & tmp_ivl_15014;
  LPM_q_ivl_15018 <= tmp_ivl_15020 & tmp_ivl_15015;
  tmp_ivl_15022 <= new_AGEMA_signal_3400 & n3912;
  LPM_q_ivl_15025 <= tmp_ivl_15027 & tmp_ivl_15022;
  new_AGEMA_signal_3677 <= tmp_ivl_15029(1);
  n3431 <= tmp_ivl_15029(0);
  tmp_ivl_15029 <= LPM_d0_ivl_15033(0 + 1 downto 0);
  tmp_ivl_15034 <= new_AGEMA_signal_3677 & n3431;
  LPM_q_ivl_15037 <= tmp_ivl_15039 & tmp_ivl_15034;
  tmp_ivl_15041 <= new_AGEMA_signal_2675 & n3430;
  LPM_q_ivl_15044 <= tmp_ivl_15046 & tmp_ivl_15041;
  new_AGEMA_signal_3957 <= tmp_ivl_15048(1);
  n3436 <= tmp_ivl_15048(0);
  tmp_ivl_15048 <= LPM_d0_ivl_15052(0 + 1 downto 0);
  tmp_ivl_15053 <= new_AGEMA_signal_4252 & n3432;
  LPM_q_ivl_15056 <= tmp_ivl_15058 & tmp_ivl_15053;
  tmp_ivl_15060 <= new_AGEMA_signal_3957 & n3436;
  LPM_q_ivl_15063 <= tmp_ivl_15065 & tmp_ivl_15060;
  tmp_ivl_15067 <= tmp_ivl_15071(1);
  tmp_ivl_15069 <= tmp_ivl_15071(0);
  tmp_ivl_15071 <= LPM_d0_ivl_15075(0 + 1 downto 0);
  tmp_ivl_15076 <= new_AGEMA_signal_3909 & n3433;
  LPM_q_ivl_15079 <= tmp_ivl_15081 & tmp_ivl_15076;
  tmp_ivl_15083 <= new_AGEMA_signal_3933 & n3745;
  LPM_q_ivl_15086 <= tmp_ivl_15088 & tmp_ivl_15083;
  new_AGEMA_signal_4253 <= tmp_ivl_15090(1);
  n3434 <= tmp_ivl_15090(0);
  tmp_ivl_15090 <= LPM_d0_ivl_15094(0 + 1 downto 0);
  tmp_ivl_15095 <= new_AGEMA_signal_4253 & n3434;
  LPM_q_ivl_15098 <= tmp_ivl_15100 & tmp_ivl_15095;
  tmp_ivl_15102 <= new_AGEMA_signal_3957 & n3436;
  LPM_q_ivl_15105 <= tmp_ivl_15107 & tmp_ivl_15102;
  tmp_ivl_15109 <= tmp_ivl_15113(1);
  tmp_ivl_15111 <= tmp_ivl_15113(0);
  tmp_ivl_15113 <= LPM_d0_ivl_15117(0 + 1 downto 0);
  tmp_ivl_15118 <= new_AGEMA_signal_3948 & n3884;
  LPM_q_ivl_15121 <= tmp_ivl_15123 & tmp_ivl_15118;
  tmp_ivl_15125 <= new_AGEMA_signal_3952 & n3435;
  LPM_q_ivl_15128 <= tmp_ivl_15130 & tmp_ivl_15125;
  new_AGEMA_signal_4254 <= tmp_ivl_15132(1);
  n3437 <= tmp_ivl_15132(0);
  tmp_ivl_15132 <= LPM_d0_ivl_15136(0 + 1 downto 0);
  tmp_ivl_15137 <= new_AGEMA_signal_4254 & n3437;
  LPM_q_ivl_15140 <= tmp_ivl_15142 & tmp_ivl_15137;
  tmp_ivl_15144 <= new_AGEMA_signal_3957 & n3436;
  LPM_q_ivl_15147 <= tmp_ivl_15149 & tmp_ivl_15144;
  tmp_ivl_15151 <= tmp_ivl_15155(1);
  tmp_ivl_15153 <= tmp_ivl_15155(0);
  tmp_ivl_15155 <= LPM_d0_ivl_15159(0 + 1 downto 0);
  tmp_ivl_15161 <= z0(11);
  tmp_ivl_15162 <= new_AGEMA_signal_3227 & tmp_ivl_15161;
  LPM_q_ivl_15165 <= tmp_ivl_15167 & tmp_ivl_15162;
  tmp_ivl_15170 <= state_in_s1(51);
  tmp_ivl_15172 <= state_in_s0(51);
  tmp_ivl_15173 <= tmp_ivl_15170 & tmp_ivl_15172;
  LPM_q_ivl_15176 <= tmp_ivl_15178 & tmp_ivl_15173;
  new_AGEMA_signal_3401 <= tmp_ivl_15180(1);
  n3448 <= tmp_ivl_15180(0);
  tmp_ivl_15180 <= LPM_d0_ivl_15184(0 + 1 downto 0);
  tmp_ivl_15185 <= new_AGEMA_signal_3401 & n3448;
  LPM_q_ivl_15188 <= tmp_ivl_15190 & tmp_ivl_15185;
  tmp_ivl_15192 <= new_AGEMA_signal_3307 & n3438;
  LPM_q_ivl_15195 <= tmp_ivl_15197 & tmp_ivl_15192;
  new_AGEMA_signal_3678 <= tmp_ivl_15199(1);
  n3704 <= tmp_ivl_15199(0);
  tmp_ivl_15199 <= LPM_d0_ivl_15203(0 + 1 downto 0);
  tmp_ivl_15204 <= new_AGEMA_signal_3360 & n3440;
  LPM_q_ivl_15207 <= tmp_ivl_15209 & tmp_ivl_15204;
  tmp_ivl_15211 <= new_AGEMA_signal_3315 & n3439;
  LPM_q_ivl_15214 <= tmp_ivl_15216 & tmp_ivl_15211;
  new_AGEMA_signal_3679 <= tmp_ivl_15218(1);
  n3671 <= tmp_ivl_15218(0);
  tmp_ivl_15218 <= LPM_d0_ivl_15222(0 + 1 downto 0);
  tmp_ivl_15223 <= new_AGEMA_signal_3678 & n3704;
  LPM_q_ivl_15226 <= tmp_ivl_15228 & tmp_ivl_15223;
  tmp_ivl_15230 <= new_AGEMA_signal_3679 & n3671;
  LPM_q_ivl_15233 <= tmp_ivl_15235 & tmp_ivl_15230;
  new_AGEMA_signal_3958 <= tmp_ivl_15237(1);
  n3443 <= tmp_ivl_15237(0);
  tmp_ivl_15237 <= LPM_d0_ivl_15241(0 + 1 downto 0);
  tmp_ivl_15242 <= new_AGEMA_signal_3341 & n3442;
  LPM_q_ivl_15245 <= tmp_ivl_15247 & tmp_ivl_15242;
  tmp_ivl_15249 <= new_AGEMA_signal_3297 & n3441;
  LPM_q_ivl_15252 <= tmp_ivl_15254 & tmp_ivl_15249;
  new_AGEMA_signal_3680 <= tmp_ivl_15256(1);
  n3667 <= tmp_ivl_15256(0);
  tmp_ivl_15256 <= LPM_d0_ivl_15260(0 + 1 downto 0);
  tmp_ivl_15261 <= new_AGEMA_signal_3958 & n3443;
  LPM_q_ivl_15264 <= tmp_ivl_15266 & tmp_ivl_15261;
  tmp_ivl_15268 <= new_AGEMA_signal_3680 & n3667;
  LPM_q_ivl_15271 <= tmp_ivl_15273 & tmp_ivl_15268;
  tmp_ivl_15275 <= tmp_ivl_15279(1);
  tmp_ivl_15277 <= tmp_ivl_15279(0);
  tmp_ivl_15279 <= LPM_d0_ivl_15283(0 + 1 downto 0);
  tmp_ivl_15285 <= z1(36);
  tmp_ivl_15286 <= new_AGEMA_signal_3017 & tmp_ivl_15285;
  LPM_q_ivl_15289 <= tmp_ivl_15291 & tmp_ivl_15286;
  tmp_ivl_15294 <= state_in_s1(284);
  tmp_ivl_15296 <= state_in_s0(284);
  tmp_ivl_15297 <= tmp_ivl_15294 & tmp_ivl_15296;
  LPM_q_ivl_15300 <= tmp_ivl_15302 & tmp_ivl_15297;
  new_AGEMA_signal_3402 <= tmp_ivl_15304(1);
  n3446 <= tmp_ivl_15304(0);
  tmp_ivl_15304 <= LPM_d0_ivl_15308(0 + 1 downto 0);
  tmp_ivl_15310 <= state_in_s1(92);
  tmp_ivl_15312 <= state_in_s0(92);
  tmp_ivl_15313 <= tmp_ivl_15310 & tmp_ivl_15312;
  LPM_q_ivl_15316 <= tmp_ivl_15318 & tmp_ivl_15313;
  tmp_ivl_15320 <= new_AGEMA_signal_3396 & n3444;
  LPM_q_ivl_15323 <= tmp_ivl_15325 & tmp_ivl_15320;
  new_AGEMA_signal_3681 <= tmp_ivl_15327(1);
  n3445 <= tmp_ivl_15327(0);
  tmp_ivl_15327 <= LPM_d0_ivl_15331(0 + 1 downto 0);
  tmp_ivl_15332 <= new_AGEMA_signal_3402 & n3446;
  LPM_q_ivl_15335 <= tmp_ivl_15337 & tmp_ivl_15332;
  tmp_ivl_15339 <= new_AGEMA_signal_3681 & n3445;
  LPM_q_ivl_15342 <= tmp_ivl_15344 & tmp_ivl_15339;
  new_AGEMA_signal_3959 <= tmp_ivl_15346(1);
  n3541 <= tmp_ivl_15346(0);
  tmp_ivl_15346 <= LPM_d0_ivl_15350(0 + 1 downto 0);
  tmp_ivl_15351 <= new_AGEMA_signal_3908 & n3447;
  LPM_q_ivl_15354 <= tmp_ivl_15356 & tmp_ivl_15351;
  tmp_ivl_15358 <= new_AGEMA_signal_3959 & n3541;
  LPM_q_ivl_15361 <= tmp_ivl_15363 & tmp_ivl_15358;
  new_AGEMA_signal_4256 <= tmp_ivl_15365(1);
  n3451 <= tmp_ivl_15365(0);
  tmp_ivl_15365 <= LPM_d0_ivl_15369(0 + 1 downto 0);
  tmp_ivl_15371 <= z1(11);
  tmp_ivl_15372 <= new_AGEMA_signal_2992 & tmp_ivl_15371;
  LPM_q_ivl_15375 <= tmp_ivl_15377 & tmp_ivl_15372;
  tmp_ivl_15379 <= new_AGEMA_signal_3401 & n3448;
  LPM_q_ivl_15382 <= tmp_ivl_15384 & tmp_ivl_15379;
  new_AGEMA_signal_3682 <= tmp_ivl_15386(1);
  n3450 <= tmp_ivl_15386(0);
  tmp_ivl_15386 <= LPM_d0_ivl_15390(0 + 1 downto 0);
  tmp_ivl_15391 <= new_AGEMA_signal_3682 & n3450;
  LPM_q_ivl_15394 <= tmp_ivl_15396 & tmp_ivl_15391;
  tmp_ivl_15398 <= new_AGEMA_signal_2677 & n3449;
  LPM_q_ivl_15401 <= tmp_ivl_15403 & tmp_ivl_15398;
  new_AGEMA_signal_3960 <= tmp_ivl_15405(1);
  n3472 <= tmp_ivl_15405(0);
  tmp_ivl_15405 <= LPM_d0_ivl_15409(0 + 1 downto 0);
  tmp_ivl_15410 <= new_AGEMA_signal_4256 & n3451;
  LPM_q_ivl_15413 <= tmp_ivl_15415 & tmp_ivl_15410;
  tmp_ivl_15417 <= new_AGEMA_signal_3960 & n3472;
  LPM_q_ivl_15420 <= tmp_ivl_15422 & tmp_ivl_15417;
  tmp_ivl_15424 <= tmp_ivl_15428(1);
  tmp_ivl_15426 <= tmp_ivl_15428(0);
  tmp_ivl_15428 <= LPM_d0_ivl_15432(0 + 1 downto 0);
  tmp_ivl_15433 <= new_AGEMA_signal_3932 & n3751;
  LPM_q_ivl_15436 <= tmp_ivl_15438 & tmp_ivl_15433;
  tmp_ivl_15440 <= new_AGEMA_signal_3936 & n3468;
  LPM_q_ivl_15443 <= tmp_ivl_15445 & tmp_ivl_15440;
  new_AGEMA_signal_4257 <= tmp_ivl_15447(1);
  n3452 <= tmp_ivl_15447(0);
  tmp_ivl_15447 <= LPM_d0_ivl_15451(0 + 1 downto 0);
  tmp_ivl_15452 <= new_AGEMA_signal_4257 & n3452;
  LPM_q_ivl_15455 <= tmp_ivl_15457 & tmp_ivl_15452;
  tmp_ivl_15459 <= new_AGEMA_signal_3960 & n3472;
  LPM_q_ivl_15462 <= tmp_ivl_15464 & tmp_ivl_15459;
  tmp_ivl_15466 <= tmp_ivl_15470(1);
  tmp_ivl_15468 <= tmp_ivl_15470(0);
  tmp_ivl_15470 <= LPM_d0_ivl_15474(0 + 1 downto 0);
  tmp_ivl_15475 <= new_AGEMA_signal_3599 & n3454;
  LPM_q_ivl_15478 <= tmp_ivl_15480 & tmp_ivl_15475;
  tmp_ivl_15482 <= new_AGEMA_signal_3628 & n3453;
  LPM_q_ivl_15485 <= tmp_ivl_15487 & tmp_ivl_15482;
  new_AGEMA_signal_3961 <= tmp_ivl_15489(1);
  n3455 <= tmp_ivl_15489(0);
  tmp_ivl_15489 <= LPM_d0_ivl_15493(0 + 1 downto 0);
  tmp_ivl_15495 <= state_in_s1(197);
  tmp_ivl_15497 <= state_in_s0(197);
  tmp_ivl_15498 <= tmp_ivl_15495 & tmp_ivl_15497;
  LPM_q_ivl_15501 <= tmp_ivl_15503 & tmp_ivl_15498;
  tmp_ivl_15506 <= z4(61);
  tmp_ivl_15507 <= new_AGEMA_signal_3168 & tmp_ivl_15506;
  LPM_q_ivl_15510 <= tmp_ivl_15512 & tmp_ivl_15507;
  new_AGEMA_signal_3403 <= tmp_ivl_15514(1);
  n3680 <= tmp_ivl_15514(0);
  tmp_ivl_15514 <= LPM_d0_ivl_15518(0 + 1 downto 0);
  tmp_ivl_15520 <= state_in_s1(261);
  tmp_ivl_15522 <= state_in_s0(261);
  tmp_ivl_15523 <= tmp_ivl_15520 & tmp_ivl_15522;
  LPM_q_ivl_15526 <= tmp_ivl_15528 & tmp_ivl_15523;
  tmp_ivl_15530 <= new_AGEMA_signal_3403 & n3680;
  LPM_q_ivl_15533 <= tmp_ivl_15535 & tmp_ivl_15530;
  new_AGEMA_signal_3683 <= tmp_ivl_15537(1);
  n3459 <= tmp_ivl_15537(0);
  tmp_ivl_15537 <= LPM_d0_ivl_15541(0 + 1 downto 0);
  tmp_ivl_15542 <= new_AGEMA_signal_3961 & n3455;
  LPM_q_ivl_15545 <= tmp_ivl_15547 & tmp_ivl_15542;
  tmp_ivl_15549 <= new_AGEMA_signal_3683 & n3459;
  LPM_q_ivl_15552 <= tmp_ivl_15554 & tmp_ivl_15549;
  tmp_ivl_15556 <= tmp_ivl_15560(1);
  tmp_ivl_15558 <= tmp_ivl_15560(0);
  tmp_ivl_15560 <= LPM_d0_ivl_15564(0 + 1 downto 0);
  tmp_ivl_15565 <= new_AGEMA_signal_3606 & n3457;
  LPM_q_ivl_15568 <= tmp_ivl_15570 & tmp_ivl_15565;
  tmp_ivl_15572 <= new_AGEMA_signal_3629 & n3456;
  LPM_q_ivl_15575 <= tmp_ivl_15577 & tmp_ivl_15572;
  new_AGEMA_signal_3962 <= tmp_ivl_15579(1);
  n3458 <= tmp_ivl_15579(0);
  tmp_ivl_15579 <= LPM_d0_ivl_15583(0 + 1 downto 0);
  tmp_ivl_15584 <= new_AGEMA_signal_3962 & n3458;
  LPM_q_ivl_15587 <= tmp_ivl_15589 & tmp_ivl_15584;
  tmp_ivl_15591 <= new_AGEMA_signal_3683 & n3459;
  LPM_q_ivl_15594 <= tmp_ivl_15596 & tmp_ivl_15591;
  tmp_ivl_15598 <= tmp_ivl_15602(1);
  tmp_ivl_15600 <= tmp_ivl_15602(0);
  tmp_ivl_15602 <= LPM_d0_ivl_15606(0 + 1 downto 0);
  tmp_ivl_15607 <= new_AGEMA_signal_3605 & n3729;
  LPM_q_ivl_15610 <= tmp_ivl_15612 & tmp_ivl_15607;
  tmp_ivl_15614 <= new_AGEMA_signal_3674 & n3725;
  LPM_q_ivl_15617 <= tmp_ivl_15619 & tmp_ivl_15614;
  new_AGEMA_signal_3963 <= tmp_ivl_15621(1);
  n3460 <= tmp_ivl_15621(0);
  tmp_ivl_15621 <= LPM_d0_ivl_15625(0 + 1 downto 0);
  tmp_ivl_15626 <= new_AGEMA_signal_3963 & n3460;
  LPM_q_ivl_15629 <= tmp_ivl_15631 & tmp_ivl_15626;
  tmp_ivl_15633 <= new_AGEMA_signal_3683 & n3459;
  LPM_q_ivl_15636 <= tmp_ivl_15638 & tmp_ivl_15633;
  tmp_ivl_15640 <= tmp_ivl_15644(1);
  tmp_ivl_15642 <= tmp_ivl_15644(0);
  tmp_ivl_15644 <= LPM_d0_ivl_15648(0 + 1 downto 0);
  tmp_ivl_15649 <= new_AGEMA_signal_3912 & n3464;
  LPM_q_ivl_15652 <= tmp_ivl_15654 & tmp_ivl_15649;
  tmp_ivl_15656 <= new_AGEMA_signal_3926 & n3617;
  LPM_q_ivl_15659 <= tmp_ivl_15661 & tmp_ivl_15656;
  new_AGEMA_signal_4261 <= tmp_ivl_15663(1);
  n3463 <= tmp_ivl_15663(0);
  tmp_ivl_15663 <= LPM_d0_ivl_15667(0 + 1 downto 0);
  tmp_ivl_15669 <= z1(14);
  tmp_ivl_15670 <= new_AGEMA_signal_2995 & tmp_ivl_15669;
  LPM_q_ivl_15673 <= tmp_ivl_15675 & tmp_ivl_15670;
  tmp_ivl_15678 <= state_in_s1(310);
  tmp_ivl_15680 <= state_in_s0(310);
  tmp_ivl_15681 <= tmp_ivl_15678 & tmp_ivl_15680;
  LPM_q_ivl_15684 <= tmp_ivl_15686 & tmp_ivl_15681;
  new_AGEMA_signal_3404 <= tmp_ivl_15688(1);
  n3462 <= tmp_ivl_15688(0);
  tmp_ivl_15688 <= LPM_d0_ivl_15692(0 + 1 downto 0);
  tmp_ivl_15694 <= z0(14);
  tmp_ivl_15695 <= new_AGEMA_signal_3228 & tmp_ivl_15694;
  LPM_q_ivl_15698 <= tmp_ivl_15700 & tmp_ivl_15695;
  tmp_ivl_15703 <= state_in_s1(54);
  tmp_ivl_15705 <= state_in_s0(54);
  tmp_ivl_15706 <= tmp_ivl_15703 & tmp_ivl_15705;
  LPM_q_ivl_15709 <= tmp_ivl_15711 & tmp_ivl_15706;
  new_AGEMA_signal_3405 <= tmp_ivl_15713(1);
  n3599 <= tmp_ivl_15713(0);
  tmp_ivl_15713 <= LPM_d0_ivl_15717(0 + 1 downto 0);
  tmp_ivl_15719 <= state_in_s1(118);
  tmp_ivl_15721 <= state_in_s0(118);
  tmp_ivl_15722 <= tmp_ivl_15719 & tmp_ivl_15721;
  LPM_q_ivl_15725 <= tmp_ivl_15727 & tmp_ivl_15722;
  tmp_ivl_15729 <= new_AGEMA_signal_3405 & n3599;
  LPM_q_ivl_15732 <= tmp_ivl_15734 & tmp_ivl_15729;
  new_AGEMA_signal_3684 <= tmp_ivl_15736(1);
  n3461 <= tmp_ivl_15736(0);
  tmp_ivl_15736 <= LPM_d0_ivl_15740(0 + 1 downto 0);
  tmp_ivl_15741 <= new_AGEMA_signal_3404 & n3462;
  LPM_q_ivl_15744 <= tmp_ivl_15746 & tmp_ivl_15741;
  tmp_ivl_15748 <= new_AGEMA_signal_3684 & n3461;
  LPM_q_ivl_15751 <= tmp_ivl_15753 & tmp_ivl_15748;
  new_AGEMA_signal_3964 <= tmp_ivl_15755(1);
  n3530 <= tmp_ivl_15755(0);
  tmp_ivl_15755 <= LPM_d0_ivl_15759(0 + 1 downto 0);
  tmp_ivl_15760 <= new_AGEMA_signal_4261 & n3463;
  LPM_q_ivl_15763 <= tmp_ivl_15765 & tmp_ivl_15760;
  tmp_ivl_15767 <= new_AGEMA_signal_3964 & n3530;
  LPM_q_ivl_15770 <= tmp_ivl_15772 & tmp_ivl_15767;
  tmp_ivl_15774 <= tmp_ivl_15778(1);
  tmp_ivl_15776 <= tmp_ivl_15778(0);
  tmp_ivl_15778 <= LPM_d0_ivl_15782(0 + 1 downto 0);
  tmp_ivl_15783 <= new_AGEMA_signal_3912 & n3464;
  LPM_q_ivl_15786 <= tmp_ivl_15788 & tmp_ivl_15783;
  tmp_ivl_15790 <= new_AGEMA_signal_3941 & n3762;
  LPM_q_ivl_15793 <= tmp_ivl_15795 & tmp_ivl_15790;
  new_AGEMA_signal_4262 <= tmp_ivl_15797(1);
  n3467 <= tmp_ivl_15797(0);
  tmp_ivl_15797 <= LPM_d0_ivl_15801(0 + 1 downto 0);
  tmp_ivl_15803 <= z1(53);
  tmp_ivl_15804 <= new_AGEMA_signal_3034 & tmp_ivl_15803;
  LPM_q_ivl_15807 <= tmp_ivl_15809 & tmp_ivl_15804;
  tmp_ivl_15812 <= state_in_s1(269);
  tmp_ivl_15814 <= state_in_s0(269);
  tmp_ivl_15815 <= tmp_ivl_15812 & tmp_ivl_15814;
  LPM_q_ivl_15818 <= tmp_ivl_15820 & tmp_ivl_15815;
  new_AGEMA_signal_3406 <= tmp_ivl_15822(1);
  n3466 <= tmp_ivl_15822(0);
  tmp_ivl_15822 <= LPM_d0_ivl_15826(0 + 1 downto 0);
  tmp_ivl_15828 <= z0(53);
  tmp_ivl_15829 <= new_AGEMA_signal_3229 & tmp_ivl_15828;
  LPM_q_ivl_15832 <= tmp_ivl_15834 & tmp_ivl_15829;
  tmp_ivl_15837 <= state_in_s1(13);
  tmp_ivl_15839 <= state_in_s0(13);
  tmp_ivl_15840 <= tmp_ivl_15837 & tmp_ivl_15839;
  LPM_q_ivl_15843 <= tmp_ivl_15845 & tmp_ivl_15840;
  new_AGEMA_signal_3407 <= tmp_ivl_15847(1);
  n3567 <= tmp_ivl_15847(0);
  tmp_ivl_15847 <= LPM_d0_ivl_15851(0 + 1 downto 0);
  tmp_ivl_15853 <= state_in_s1(77);
  tmp_ivl_15855 <= state_in_s0(77);
  tmp_ivl_15856 <= tmp_ivl_15853 & tmp_ivl_15855;
  LPM_q_ivl_15859 <= tmp_ivl_15861 & tmp_ivl_15856;
  tmp_ivl_15863 <= new_AGEMA_signal_3407 & n3567;
  LPM_q_ivl_15866 <= tmp_ivl_15868 & tmp_ivl_15863;
  new_AGEMA_signal_3685 <= tmp_ivl_15870(1);
  n3465 <= tmp_ivl_15870(0);
  tmp_ivl_15870 <= LPM_d0_ivl_15874(0 + 1 downto 0);
  tmp_ivl_15875 <= new_AGEMA_signal_3406 & n3466;
  LPM_q_ivl_15878 <= tmp_ivl_15880 & tmp_ivl_15875;
  tmp_ivl_15882 <= new_AGEMA_signal_3685 & n3465;
  LPM_q_ivl_15885 <= tmp_ivl_15887 & tmp_ivl_15882;
  new_AGEMA_signal_3965 <= tmp_ivl_15889(1);
  n3473 <= tmp_ivl_15889(0);
  tmp_ivl_15889 <= LPM_d0_ivl_15893(0 + 1 downto 0);
  tmp_ivl_15894 <= new_AGEMA_signal_4262 & n3467;
  LPM_q_ivl_15897 <= tmp_ivl_15899 & tmp_ivl_15894;
  tmp_ivl_15901 <= new_AGEMA_signal_3965 & n3473;
  LPM_q_ivl_15904 <= tmp_ivl_15906 & tmp_ivl_15901;
  tmp_ivl_15908 <= tmp_ivl_15912(1);
  tmp_ivl_15910 <= tmp_ivl_15912(0);
  tmp_ivl_15912 <= LPM_d0_ivl_15916(0 + 1 downto 0);
  tmp_ivl_15917 <= new_AGEMA_signal_3936 & n3468;
  LPM_q_ivl_15920 <= tmp_ivl_15922 & tmp_ivl_15917;
  tmp_ivl_15924 <= new_AGEMA_signal_3965 & n3473;
  LPM_q_ivl_15927 <= tmp_ivl_15929 & tmp_ivl_15924;
  new_AGEMA_signal_4263 <= tmp_ivl_15931(1);
  n3471 <= tmp_ivl_15931(0);
  tmp_ivl_15931 <= LPM_d0_ivl_15935(0 + 1 downto 0);
  tmp_ivl_15937 <= z0(28);
  tmp_ivl_15938 <= new_AGEMA_signal_3255 & tmp_ivl_15937;
  LPM_q_ivl_15941 <= tmp_ivl_15943 & tmp_ivl_15938;
  tmp_ivl_15946 <= state_in_s1(36);
  tmp_ivl_15948 <= state_in_s0(36);
  tmp_ivl_15949 <= tmp_ivl_15946 & tmp_ivl_15948;
  LPM_q_ivl_15952 <= tmp_ivl_15954 & tmp_ivl_15949;
  new_AGEMA_signal_3408 <= tmp_ivl_15956(1);
  n3475 <= tmp_ivl_15956(0);
  tmp_ivl_15956 <= LPM_d0_ivl_15960(0 + 1 downto 0);
  tmp_ivl_15962 <= z1(28);
  tmp_ivl_15963 <= new_AGEMA_signal_3009 & tmp_ivl_15962;
  LPM_q_ivl_15966 <= tmp_ivl_15968 & tmp_ivl_15963;
  tmp_ivl_15970 <= new_AGEMA_signal_3408 & n3475;
  LPM_q_ivl_15973 <= tmp_ivl_15975 & tmp_ivl_15970;
  new_AGEMA_signal_3686 <= tmp_ivl_15977(1);
  n3470 <= tmp_ivl_15977(0);
  tmp_ivl_15977 <= LPM_d0_ivl_15981(0 + 1 downto 0);
  tmp_ivl_15982 <= new_AGEMA_signal_3686 & n3470;
  LPM_q_ivl_15985 <= tmp_ivl_15987 & tmp_ivl_15982;
  tmp_ivl_15989 <= new_AGEMA_signal_2679 & n3469;
  LPM_q_ivl_15992 <= tmp_ivl_15994 & tmp_ivl_15989;
  new_AGEMA_signal_3966 <= tmp_ivl_15996(1);
  n3809 <= tmp_ivl_15996(0);
  tmp_ivl_15996 <= LPM_d0_ivl_16000(0 + 1 downto 0);
  tmp_ivl_16001 <= new_AGEMA_signal_4263 & n3471;
  LPM_q_ivl_16004 <= tmp_ivl_16006 & tmp_ivl_16001;
  tmp_ivl_16008 <= new_AGEMA_signal_3966 & n3809;
  LPM_q_ivl_16011 <= tmp_ivl_16013 & tmp_ivl_16008;
  tmp_ivl_16015 <= tmp_ivl_16019(1);
  tmp_ivl_16017 <= tmp_ivl_16019(0);
  tmp_ivl_16019 <= LPM_d0_ivl_16023(0 + 1 downto 0);
  tmp_ivl_16024 <= new_AGEMA_signal_3960 & n3472;
  LPM_q_ivl_16027 <= tmp_ivl_16029 & tmp_ivl_16024;
  tmp_ivl_16031 <= new_AGEMA_signal_3964 & n3530;
  LPM_q_ivl_16034 <= tmp_ivl_16036 & tmp_ivl_16031;
  new_AGEMA_signal_4264 <= tmp_ivl_16038(1);
  n3474 <= tmp_ivl_16038(0);
  tmp_ivl_16038 <= LPM_d0_ivl_16042(0 + 1 downto 0);
  tmp_ivl_16043 <= new_AGEMA_signal_4264 & n3474;
  LPM_q_ivl_16046 <= tmp_ivl_16048 & tmp_ivl_16043;
  tmp_ivl_16050 <= new_AGEMA_signal_3965 & n3473;
  LPM_q_ivl_16053 <= tmp_ivl_16055 & tmp_ivl_16050;
  tmp_ivl_16057 <= tmp_ivl_16061(1);
  tmp_ivl_16059 <= tmp_ivl_16061(0);
  tmp_ivl_16061 <= LPM_d0_ivl_16065(0 + 1 downto 0);
  tmp_ivl_16066 <= new_AGEMA_signal_3644 & n3705;
  LPM_q_ivl_16069 <= tmp_ivl_16071 & tmp_ivl_16066;
  tmp_ivl_16073 <= new_AGEMA_signal_3680 & n3667;
  LPM_q_ivl_16076 <= tmp_ivl_16078 & tmp_ivl_16073;
  new_AGEMA_signal_3967 <= tmp_ivl_16080(1);
  n3476 <= tmp_ivl_16080(0);
  tmp_ivl_16080 <= LPM_d0_ivl_16084(0 + 1 downto 0);
  tmp_ivl_16086 <= state_in_s1(228);
  tmp_ivl_16088 <= state_in_s0(228);
  tmp_ivl_16089 <= tmp_ivl_16086 & tmp_ivl_16088;
  LPM_q_ivl_16092 <= tmp_ivl_16094 & tmp_ivl_16089;
  tmp_ivl_16097 <= z4(28);
  tmp_ivl_16098 <= new_AGEMA_signal_3131 & tmp_ivl_16097;
  LPM_q_ivl_16101 <= tmp_ivl_16103 & tmp_ivl_16098;
  new_AGEMA_signal_3409 <= tmp_ivl_16105(1);
  n3482 <= tmp_ivl_16105(0);
  tmp_ivl_16105 <= LPM_d0_ivl_16109(0 + 1 downto 0);
  tmp_ivl_16110 <= new_AGEMA_signal_3408 & n3475;
  LPM_q_ivl_16113 <= tmp_ivl_16115 & tmp_ivl_16110;
  tmp_ivl_16117 <= new_AGEMA_signal_3409 & n3482;
  LPM_q_ivl_16120 <= tmp_ivl_16122 & tmp_ivl_16117;
  new_AGEMA_signal_3687 <= tmp_ivl_16124(1);
  n3636 <= tmp_ivl_16124(0);
  tmp_ivl_16124 <= LPM_d0_ivl_16128(0 + 1 downto 0);
  tmp_ivl_16129 <= new_AGEMA_signal_3967 & n3476;
  LPM_q_ivl_16132 <= tmp_ivl_16134 & tmp_ivl_16129;
  tmp_ivl_16136 <= new_AGEMA_signal_3687 & n3636;
  LPM_q_ivl_16139 <= tmp_ivl_16141 & tmp_ivl_16136;
  tmp_ivl_16143 <= tmp_ivl_16147(1);
  tmp_ivl_16145 <= tmp_ivl_16147(0);
  tmp_ivl_16147 <= LPM_d0_ivl_16151(0 + 1 downto 0);
  tmp_ivl_16153 <= z0(37);
  tmp_ivl_16154 <= new_AGEMA_signal_3266 & tmp_ivl_16153;
  LPM_q_ivl_16157 <= tmp_ivl_16159 & tmp_ivl_16154;
  tmp_ivl_16162 <= state_in_s1(29);
  tmp_ivl_16164 <= state_in_s0(29);
  tmp_ivl_16165 <= tmp_ivl_16162 & tmp_ivl_16164;
  LPM_q_ivl_16168 <= tmp_ivl_16170 & tmp_ivl_16165;
  new_AGEMA_signal_3410 <= tmp_ivl_16172(1);
  n3499 <= tmp_ivl_16172(0);
  tmp_ivl_16172 <= LPM_d0_ivl_16176(0 + 1 downto 0);
  tmp_ivl_16177 <= new_AGEMA_signal_3410 & n3499;
  LPM_q_ivl_16180 <= tmp_ivl_16182 & tmp_ivl_16177;
  tmp_ivl_16184 <= new_AGEMA_signal_3328 & n3477;
  LPM_q_ivl_16187 <= tmp_ivl_16189 & tmp_ivl_16184;
  new_AGEMA_signal_3688 <= tmp_ivl_16191(1);
  n3863 <= tmp_ivl_16191(0);
  tmp_ivl_16191 <= LPM_d0_ivl_16195(0 + 1 downto 0);
  tmp_ivl_16196 <= new_AGEMA_signal_3687 & n3636;
  LPM_q_ivl_16199 <= tmp_ivl_16201 & tmp_ivl_16196;
  tmp_ivl_16203 <= new_AGEMA_signal_3688 & n3863;
  LPM_q_ivl_16206 <= tmp_ivl_16208 & tmp_ivl_16203;
  new_AGEMA_signal_3968 <= tmp_ivl_16210(1);
  n3480 <= tmp_ivl_16210(0);
  tmp_ivl_16210 <= LPM_d0_ivl_16214(0 + 1 downto 0);
  tmp_ivl_16215 <= new_AGEMA_signal_3378 & n3479;
  LPM_q_ivl_16218 <= tmp_ivl_16220 & tmp_ivl_16215;
  tmp_ivl_16222 <= new_AGEMA_signal_3301 & n3478;
  LPM_q_ivl_16225 <= tmp_ivl_16227 & tmp_ivl_16222;
  new_AGEMA_signal_3689 <= tmp_ivl_16229(1);
  n3860 <= tmp_ivl_16229(0);
  tmp_ivl_16229 <= LPM_d0_ivl_16233(0 + 1 downto 0);
  tmp_ivl_16234 <= new_AGEMA_signal_3968 & n3480;
  LPM_q_ivl_16237 <= tmp_ivl_16239 & tmp_ivl_16234;
  tmp_ivl_16241 <= new_AGEMA_signal_3689 & n3860;
  LPM_q_ivl_16244 <= tmp_ivl_16246 & tmp_ivl_16241;
  tmp_ivl_16248 <= tmp_ivl_16252(1);
  tmp_ivl_16250 <= tmp_ivl_16252(0);
  tmp_ivl_16252 <= LPM_d0_ivl_16256(0 + 1 downto 0);
  tmp_ivl_16257 <= new_AGEMA_signal_3604 & n3508;
  LPM_q_ivl_16260 <= tmp_ivl_16262 & tmp_ivl_16257;
  tmp_ivl_16264 <= new_AGEMA_signal_3616 & n3481;
  LPM_q_ivl_16267 <= tmp_ivl_16269 & tmp_ivl_16264;
  new_AGEMA_signal_3969 <= tmp_ivl_16271(1);
  n3483 <= tmp_ivl_16271(0);
  tmp_ivl_16271 <= LPM_d0_ivl_16275(0 + 1 downto 0);
  tmp_ivl_16277 <= state_in_s1(292);
  tmp_ivl_16279 <= state_in_s0(292);
  tmp_ivl_16280 <= tmp_ivl_16277 & tmp_ivl_16279;
  LPM_q_ivl_16283 <= tmp_ivl_16285 & tmp_ivl_16280;
  tmp_ivl_16287 <= new_AGEMA_signal_3409 & n3482;
  LPM_q_ivl_16290 <= tmp_ivl_16292 & tmp_ivl_16287;
  new_AGEMA_signal_3690 <= tmp_ivl_16294(1);
  n3831 <= tmp_ivl_16294(0);
  tmp_ivl_16294 <= LPM_d0_ivl_16298(0 + 1 downto 0);
  tmp_ivl_16299 <= new_AGEMA_signal_3969 & n3483;
  LPM_q_ivl_16302 <= tmp_ivl_16304 & tmp_ivl_16299;
  tmp_ivl_16306 <= new_AGEMA_signal_3690 & n3831;
  LPM_q_ivl_16309 <= tmp_ivl_16311 & tmp_ivl_16306;
  tmp_ivl_16313 <= tmp_ivl_16317(1);
  tmp_ivl_16315 <= tmp_ivl_16317(0);
  tmp_ivl_16317 <= LPM_d0_ivl_16321(0 + 1 downto 0);
  tmp_ivl_16323 <= z0(24);
  tmp_ivl_16324 <= new_AGEMA_signal_3261 & tmp_ivl_16323;
  LPM_q_ivl_16327 <= tmp_ivl_16329 & tmp_ivl_16324;
  tmp_ivl_16332 <= state_in_s1(32);
  tmp_ivl_16334 <= state_in_s0(32);
  tmp_ivl_16335 <= tmp_ivl_16332 & tmp_ivl_16334;
  LPM_q_ivl_16338 <= tmp_ivl_16340 & tmp_ivl_16335;
  new_AGEMA_signal_3411 <= tmp_ivl_16342(1);
  n3591 <= tmp_ivl_16342(0);
  tmp_ivl_16342 <= LPM_d0_ivl_16346(0 + 1 downto 0);
  tmp_ivl_16347 <= new_AGEMA_signal_3411 & n3591;
  LPM_q_ivl_16350 <= tmp_ivl_16352 & tmp_ivl_16347;
  tmp_ivl_16354 <= new_AGEMA_signal_3358 & n3484;
  LPM_q_ivl_16357 <= tmp_ivl_16359 & tmp_ivl_16354;
  new_AGEMA_signal_3691 <= tmp_ivl_16361(1);
  n3918 <= tmp_ivl_16361(0);
  tmp_ivl_16361 <= LPM_d0_ivl_16365(0 + 1 downto 0);
  tmp_ivl_16366 <= new_AGEMA_signal_3347 & n3486;
  LPM_q_ivl_16369 <= tmp_ivl_16371 & tmp_ivl_16366;
  tmp_ivl_16373 <= new_AGEMA_signal_3385 & n3485;
  LPM_q_ivl_16376 <= tmp_ivl_16378 & tmp_ivl_16373;
  new_AGEMA_signal_3692 <= tmp_ivl_16380(1);
  n3826 <= tmp_ivl_16380(0);
  tmp_ivl_16380 <= LPM_d0_ivl_16384(0 + 1 downto 0);
  tmp_ivl_16385 <= new_AGEMA_signal_3691 & n3918;
  LPM_q_ivl_16388 <= tmp_ivl_16390 & tmp_ivl_16385;
  tmp_ivl_16392 <= new_AGEMA_signal_3692 & n3826;
  LPM_q_ivl_16395 <= tmp_ivl_16397 & tmp_ivl_16392;
  new_AGEMA_signal_3970 <= tmp_ivl_16399(1);
  n3488 <= tmp_ivl_16399(0);
  tmp_ivl_16399 <= LPM_d0_ivl_16403(0 + 1 downto 0);
  tmp_ivl_16405 <= z0(15);
  tmp_ivl_16406 <= new_AGEMA_signal_3224 & tmp_ivl_16405;
  LPM_q_ivl_16409 <= tmp_ivl_16411 & tmp_ivl_16406;
  tmp_ivl_16414 <= state_in_s1(55);
  tmp_ivl_16416 <= state_in_s0(55);
  tmp_ivl_16417 <= tmp_ivl_16414 & tmp_ivl_16416;
  LPM_q_ivl_16420 <= tmp_ivl_16422 & tmp_ivl_16417;
  new_AGEMA_signal_3412 <= tmp_ivl_16424(1);
  n3489 <= tmp_ivl_16424(0);
  tmp_ivl_16424 <= LPM_d0_ivl_16428(0 + 1 downto 0);
  tmp_ivl_16429 <= new_AGEMA_signal_3412 & n3489;
  LPM_q_ivl_16432 <= tmp_ivl_16434 & tmp_ivl_16429;
  tmp_ivl_16436 <= new_AGEMA_signal_3296 & n3487;
  LPM_q_ivl_16439 <= tmp_ivl_16441 & tmp_ivl_16436;
  new_AGEMA_signal_3693 <= tmp_ivl_16443(1);
  n3823 <= tmp_ivl_16443(0);
  tmp_ivl_16443 <= LPM_d0_ivl_16447(0 + 1 downto 0);
  tmp_ivl_16448 <= new_AGEMA_signal_3970 & n3488;
  LPM_q_ivl_16451 <= tmp_ivl_16453 & tmp_ivl_16448;
  tmp_ivl_16455 <= new_AGEMA_signal_3693 & n3823;
  LPM_q_ivl_16458 <= tmp_ivl_16460 & tmp_ivl_16455;
  tmp_ivl_16462 <= tmp_ivl_16466(1);
  tmp_ivl_16464 <= tmp_ivl_16466(0);
  tmp_ivl_16466 <= LPM_d0_ivl_16470(0 + 1 downto 0);
  tmp_ivl_16471 <= new_AGEMA_signal_3917 & n3515;
  LPM_q_ivl_16474 <= tmp_ivl_16476 & tmp_ivl_16471;
  tmp_ivl_16478 <= new_AGEMA_signal_3920 & n3648;
  LPM_q_ivl_16481 <= tmp_ivl_16483 & tmp_ivl_16478;
  new_AGEMA_signal_4269 <= tmp_ivl_16485(1);
  n3492 <= tmp_ivl_16485(0);
  tmp_ivl_16485 <= LPM_d0_ivl_16489(0 + 1 downto 0);
  tmp_ivl_16491 <= z1(15);
  tmp_ivl_16492 <= new_AGEMA_signal_2996 & tmp_ivl_16491;
  LPM_q_ivl_16495 <= tmp_ivl_16497 & tmp_ivl_16492;
  tmp_ivl_16500 <= state_in_s1(311);
  tmp_ivl_16502 <= state_in_s0(311);
  tmp_ivl_16503 <= tmp_ivl_16500 & tmp_ivl_16502;
  LPM_q_ivl_16506 <= tmp_ivl_16508 & tmp_ivl_16503;
  new_AGEMA_signal_3413 <= tmp_ivl_16510(1);
  n3491 <= tmp_ivl_16510(0);
  tmp_ivl_16510 <= LPM_d0_ivl_16514(0 + 1 downto 0);
  tmp_ivl_16516 <= state_in_s1(119);
  tmp_ivl_16518 <= state_in_s0(119);
  tmp_ivl_16519 <= tmp_ivl_16516 & tmp_ivl_16518;
  LPM_q_ivl_16522 <= tmp_ivl_16524 & tmp_ivl_16519;
  tmp_ivl_16526 <= new_AGEMA_signal_3412 & n3489;
  LPM_q_ivl_16529 <= tmp_ivl_16531 & tmp_ivl_16526;
  new_AGEMA_signal_3694 <= tmp_ivl_16533(1);
  n3490 <= tmp_ivl_16533(0);
  tmp_ivl_16533 <= LPM_d0_ivl_16537(0 + 1 downto 0);
  tmp_ivl_16538 <= new_AGEMA_signal_3413 & n3491;
  LPM_q_ivl_16541 <= tmp_ivl_16543 & tmp_ivl_16538;
  tmp_ivl_16545 <= new_AGEMA_signal_3694 & n3490;
  LPM_q_ivl_16548 <= tmp_ivl_16550 & tmp_ivl_16545;
  new_AGEMA_signal_3971 <= tmp_ivl_16552(1);
  n3554 <= tmp_ivl_16552(0);
  tmp_ivl_16552 <= LPM_d0_ivl_16556(0 + 1 downto 0);
  tmp_ivl_16557 <= new_AGEMA_signal_4269 & n3492;
  LPM_q_ivl_16560 <= tmp_ivl_16562 & tmp_ivl_16557;
  tmp_ivl_16564 <= new_AGEMA_signal_3971 & n3554;
  LPM_q_ivl_16567 <= tmp_ivl_16569 & tmp_ivl_16564;
  tmp_ivl_16571 <= tmp_ivl_16575(1);
  tmp_ivl_16573 <= tmp_ivl_16575(0);
  tmp_ivl_16575 <= LPM_d0_ivl_16579(0 + 1 downto 0);
  tmp_ivl_16581 <= z0(12);
  tmp_ivl_16582 <= new_AGEMA_signal_3225 & tmp_ivl_16581;
  LPM_q_ivl_16585 <= tmp_ivl_16587 & tmp_ivl_16582;
  tmp_ivl_16590 <= state_in_s1(52);
  tmp_ivl_16592 <= state_in_s0(52);
  tmp_ivl_16593 <= tmp_ivl_16590 & tmp_ivl_16592;
  LPM_q_ivl_16596 <= tmp_ivl_16598 & tmp_ivl_16593;
  new_AGEMA_signal_3414 <= tmp_ivl_16600(1);
  n3503 <= tmp_ivl_16600(0);
  tmp_ivl_16600 <= LPM_d0_ivl_16604(0 + 1 downto 0);
  tmp_ivl_16605 <= new_AGEMA_signal_3414 & n3503;
  LPM_q_ivl_16608 <= tmp_ivl_16610 & tmp_ivl_16605;
  tmp_ivl_16612 <= new_AGEMA_signal_3312 & n3493;
  LPM_q_ivl_16615 <= tmp_ivl_16617 & tmp_ivl_16612;
  new_AGEMA_signal_3695 <= tmp_ivl_16619(1);
  n3799 <= tmp_ivl_16619(0);
  tmp_ivl_16619 <= LPM_d0_ivl_16623(0 + 1 downto 0);
  tmp_ivl_16624 <= new_AGEMA_signal_3352 & n3495;
  LPM_q_ivl_16627 <= tmp_ivl_16629 & tmp_ivl_16624;
  tmp_ivl_16631 <= new_AGEMA_signal_3330 & n3494;
  LPM_q_ivl_16634 <= tmp_ivl_16636 & tmp_ivl_16631;
  new_AGEMA_signal_3696 <= tmp_ivl_16638(1);
  n3712 <= tmp_ivl_16638(0);
  tmp_ivl_16638 <= LPM_d0_ivl_16642(0 + 1 downto 0);
  tmp_ivl_16643 <= new_AGEMA_signal_3695 & n3799;
  LPM_q_ivl_16646 <= tmp_ivl_16648 & tmp_ivl_16643;
  tmp_ivl_16650 <= new_AGEMA_signal_3696 & n3712;
  LPM_q_ivl_16653 <= tmp_ivl_16655 & tmp_ivl_16650;
  new_AGEMA_signal_3972 <= tmp_ivl_16657(1);
  n3498 <= tmp_ivl_16657(0);
  tmp_ivl_16657 <= LPM_d0_ivl_16661(0 + 1 downto 0);
  tmp_ivl_16662 <= new_AGEMA_signal_3348 & n3497;
  LPM_q_ivl_16665 <= tmp_ivl_16667 & tmp_ivl_16662;
  tmp_ivl_16669 <= new_AGEMA_signal_3344 & n3496;
  LPM_q_ivl_16672 <= tmp_ivl_16674 & tmp_ivl_16669;
  new_AGEMA_signal_3697 <= tmp_ivl_16676(1);
  n3708 <= tmp_ivl_16676(0);
  tmp_ivl_16676 <= LPM_d0_ivl_16680(0 + 1 downto 0);
  tmp_ivl_16681 <= new_AGEMA_signal_3972 & n3498;
  LPM_q_ivl_16684 <= tmp_ivl_16686 & tmp_ivl_16681;
  tmp_ivl_16688 <= new_AGEMA_signal_3697 & n3708;
  LPM_q_ivl_16691 <= tmp_ivl_16693 & tmp_ivl_16688;
  tmp_ivl_16695 <= tmp_ivl_16699(1);
  tmp_ivl_16697 <= tmp_ivl_16699(0);
  tmp_ivl_16699 <= LPM_d0_ivl_16703(0 + 1 downto 0);
  tmp_ivl_16705 <= z1(37);
  tmp_ivl_16706 <= new_AGEMA_signal_3018 & tmp_ivl_16705;
  LPM_q_ivl_16709 <= tmp_ivl_16711 & tmp_ivl_16706;
  tmp_ivl_16714 <= state_in_s1(285);
  tmp_ivl_16716 <= state_in_s0(285);
  tmp_ivl_16717 <= tmp_ivl_16714 & tmp_ivl_16716;
  LPM_q_ivl_16720 <= tmp_ivl_16722 & tmp_ivl_16717;
  new_AGEMA_signal_3415 <= tmp_ivl_16724(1);
  n3501 <= tmp_ivl_16724(0);
  tmp_ivl_16724 <= LPM_d0_ivl_16728(0 + 1 downto 0);
  tmp_ivl_16730 <= state_in_s1(93);
  tmp_ivl_16732 <= state_in_s0(93);
  tmp_ivl_16733 <= tmp_ivl_16730 & tmp_ivl_16732;
  LPM_q_ivl_16736 <= tmp_ivl_16738 & tmp_ivl_16733;
  tmp_ivl_16740 <= new_AGEMA_signal_3410 & n3499;
  LPM_q_ivl_16743 <= tmp_ivl_16745 & tmp_ivl_16740;
  new_AGEMA_signal_3698 <= tmp_ivl_16747(1);
  n3500 <= tmp_ivl_16747(0);
  tmp_ivl_16747 <= LPM_d0_ivl_16751(0 + 1 downto 0);
  tmp_ivl_16752 <= new_AGEMA_signal_3415 & n3501;
  LPM_q_ivl_16755 <= tmp_ivl_16757 & tmp_ivl_16752;
  tmp_ivl_16759 <= new_AGEMA_signal_3698 & n3500;
  LPM_q_ivl_16762 <= tmp_ivl_16764 & tmp_ivl_16759;
  new_AGEMA_signal_3973 <= tmp_ivl_16766(1);
  n3571 <= tmp_ivl_16766(0);
  tmp_ivl_16766 <= LPM_d0_ivl_16770(0 + 1 downto 0);
  tmp_ivl_16771 <= new_AGEMA_signal_3911 & n3502;
  LPM_q_ivl_16774 <= tmp_ivl_16776 & tmp_ivl_16771;
  tmp_ivl_16778 <= new_AGEMA_signal_3973 & n3571;
  LPM_q_ivl_16781 <= tmp_ivl_16783 & tmp_ivl_16778;
  new_AGEMA_signal_4271 <= tmp_ivl_16785(1);
  n3506 <= tmp_ivl_16785(0);
  tmp_ivl_16785 <= LPM_d0_ivl_16789(0 + 1 downto 0);
  tmp_ivl_16791 <= z1(12);
  tmp_ivl_16792 <= new_AGEMA_signal_2993 & tmp_ivl_16791;
  LPM_q_ivl_16795 <= tmp_ivl_16797 & tmp_ivl_16792;
  tmp_ivl_16800 <= state_in_s1(308);
  tmp_ivl_16802 <= state_in_s0(308);
  tmp_ivl_16803 <= tmp_ivl_16800 & tmp_ivl_16802;
  LPM_q_ivl_16806 <= tmp_ivl_16808 & tmp_ivl_16803;
  new_AGEMA_signal_3416 <= tmp_ivl_16810(1);
  n3505 <= tmp_ivl_16810(0);
  tmp_ivl_16810 <= LPM_d0_ivl_16814(0 + 1 downto 0);
  tmp_ivl_16816 <= state_in_s1(116);
  tmp_ivl_16818 <= state_in_s0(116);
  tmp_ivl_16819 <= tmp_ivl_16816 & tmp_ivl_16818;
  LPM_q_ivl_16822 <= tmp_ivl_16824 & tmp_ivl_16819;
  tmp_ivl_16826 <= new_AGEMA_signal_3414 & n3503;
  LPM_q_ivl_16829 <= tmp_ivl_16831 & tmp_ivl_16826;
  new_AGEMA_signal_3699 <= tmp_ivl_16833(1);
  n3504 <= tmp_ivl_16833(0);
  tmp_ivl_16833 <= LPM_d0_ivl_16837(0 + 1 downto 0);
  tmp_ivl_16838 <= new_AGEMA_signal_3416 & n3505;
  LPM_q_ivl_16841 <= tmp_ivl_16843 & tmp_ivl_16838;
  tmp_ivl_16845 <= new_AGEMA_signal_3699 & n3504;
  LPM_q_ivl_16848 <= tmp_ivl_16850 & tmp_ivl_16845;
  new_AGEMA_signal_3974 <= tmp_ivl_16852(1);
  n3523 <= tmp_ivl_16852(0);
  tmp_ivl_16852 <= LPM_d0_ivl_16856(0 + 1 downto 0);
  tmp_ivl_16857 <= new_AGEMA_signal_4271 & n3506;
  LPM_q_ivl_16860 <= tmp_ivl_16862 & tmp_ivl_16857;
  tmp_ivl_16864 <= new_AGEMA_signal_3974 & n3523;
  LPM_q_ivl_16867 <= tmp_ivl_16869 & tmp_ivl_16864;
  tmp_ivl_16871 <= tmp_ivl_16875(1);
  tmp_ivl_16873 <= tmp_ivl_16875(0);
  tmp_ivl_16875 <= LPM_d0_ivl_16879(0 + 1 downto 0);
  tmp_ivl_16880 <= new_AGEMA_signal_3940 & n3767;
  LPM_q_ivl_16883 <= tmp_ivl_16885 & tmp_ivl_16880;
  tmp_ivl_16887 <= new_AGEMA_signal_3944 & n3519;
  LPM_q_ivl_16890 <= tmp_ivl_16892 & tmp_ivl_16887;
  new_AGEMA_signal_4272 <= tmp_ivl_16894(1);
  n3507 <= tmp_ivl_16894(0);
  tmp_ivl_16894 <= LPM_d0_ivl_16898(0 + 1 downto 0);
  tmp_ivl_16899 <= new_AGEMA_signal_4272 & n3507;
  LPM_q_ivl_16902 <= tmp_ivl_16904 & tmp_ivl_16899;
  tmp_ivl_16906 <= new_AGEMA_signal_3974 & n3523;
  LPM_q_ivl_16909 <= tmp_ivl_16911 & tmp_ivl_16906;
  tmp_ivl_16913 <= tmp_ivl_16917(1);
  tmp_ivl_16915 <= tmp_ivl_16917(0);
  tmp_ivl_16917 <= LPM_d0_ivl_16921(0 + 1 downto 0);
  tmp_ivl_16922 <= new_AGEMA_signal_3604 & n3508;
  LPM_q_ivl_16925 <= tmp_ivl_16927 & tmp_ivl_16922;
  tmp_ivl_16929 <= new_AGEMA_signal_3610 & n3686;
  LPM_q_ivl_16932 <= tmp_ivl_16934 & tmp_ivl_16929;
  new_AGEMA_signal_3975 <= tmp_ivl_16936(1);
  n3509 <= tmp_ivl_16936(0);
  tmp_ivl_16936 <= LPM_d0_ivl_16940(0 + 1 downto 0);
  tmp_ivl_16942 <= state_in_s1(198);
  tmp_ivl_16944 <= state_in_s0(198);
  tmp_ivl_16945 <= tmp_ivl_16942 & tmp_ivl_16944;
  LPM_q_ivl_16948 <= tmp_ivl_16950 & tmp_ivl_16945;
  tmp_ivl_16953 <= z4(62);
  tmp_ivl_16954 <= new_AGEMA_signal_3169 & tmp_ivl_16953;
  LPM_q_ivl_16957 <= tmp_ivl_16959 & tmp_ivl_16954;
  new_AGEMA_signal_3417 <= tmp_ivl_16961(1);
  n3565 <= tmp_ivl_16961(0);
  tmp_ivl_16961 <= LPM_d0_ivl_16965(0 + 1 downto 0);
  tmp_ivl_16967 <= state_in_s1(262);
  tmp_ivl_16969 <= state_in_s0(262);
  tmp_ivl_16970 <= tmp_ivl_16967 & tmp_ivl_16969;
  LPM_q_ivl_16973 <= tmp_ivl_16975 & tmp_ivl_16970;
  tmp_ivl_16977 <= new_AGEMA_signal_3417 & n3565;
  LPM_q_ivl_16980 <= tmp_ivl_16982 & tmp_ivl_16977;
  new_AGEMA_signal_3700 <= tmp_ivl_16984(1);
  n3513 <= tmp_ivl_16984(0);
  tmp_ivl_16984 <= LPM_d0_ivl_16988(0 + 1 downto 0);
  tmp_ivl_16989 <= new_AGEMA_signal_3975 & n3509;
  LPM_q_ivl_16992 <= tmp_ivl_16994 & tmp_ivl_16989;
  tmp_ivl_16996 <= new_AGEMA_signal_3700 & n3513;
  LPM_q_ivl_16999 <= tmp_ivl_17001 & tmp_ivl_16996;
  tmp_ivl_17003 <= tmp_ivl_17007(1);
  tmp_ivl_17005 <= tmp_ivl_17007(0);
  tmp_ivl_17007 <= LPM_d0_ivl_17011(0 + 1 downto 0);
  tmp_ivl_17012 <= new_AGEMA_signal_3611 & n3511;
  LPM_q_ivl_17015 <= tmp_ivl_17017 & tmp_ivl_17012;
  tmp_ivl_17019 <= new_AGEMA_signal_3621 & n3510;
  LPM_q_ivl_17022 <= tmp_ivl_17024 & tmp_ivl_17019;
  new_AGEMA_signal_3976 <= tmp_ivl_17026(1);
  n3512 <= tmp_ivl_17026(0);
  tmp_ivl_17026 <= LPM_d0_ivl_17030(0 + 1 downto 0);
  tmp_ivl_17031 <= new_AGEMA_signal_3976 & n3512;
  LPM_q_ivl_17034 <= tmp_ivl_17036 & tmp_ivl_17031;
  tmp_ivl_17038 <= new_AGEMA_signal_3700 & n3513;
  LPM_q_ivl_17041 <= tmp_ivl_17043 & tmp_ivl_17038;
  tmp_ivl_17045 <= tmp_ivl_17049(1);
  tmp_ivl_17047 <= tmp_ivl_17049(0);
  tmp_ivl_17049 <= LPM_d0_ivl_17053(0 + 1 downto 0);
  tmp_ivl_17054 <= new_AGEMA_signal_3620 & n3835;
  LPM_q_ivl_17057 <= tmp_ivl_17059 & tmp_ivl_17054;
  tmp_ivl_17061 <= new_AGEMA_signal_3690 & n3831;
  LPM_q_ivl_17064 <= tmp_ivl_17066 & tmp_ivl_17061;
  new_AGEMA_signal_3977 <= tmp_ivl_17068(1);
  n3514 <= tmp_ivl_17068(0);
  tmp_ivl_17068 <= LPM_d0_ivl_17072(0 + 1 downto 0);
  tmp_ivl_17073 <= new_AGEMA_signal_3977 & n3514;
  LPM_q_ivl_17076 <= tmp_ivl_17078 & tmp_ivl_17073;
  tmp_ivl_17080 <= new_AGEMA_signal_3700 & n3513;
  LPM_q_ivl_17083 <= tmp_ivl_17085 & tmp_ivl_17080;
  tmp_ivl_17087 <= tmp_ivl_17091(1);
  tmp_ivl_17089 <= tmp_ivl_17091(0);
  tmp_ivl_17091 <= LPM_d0_ivl_17095(0 + 1 downto 0);
  tmp_ivl_17096 <= new_AGEMA_signal_3917 & n3515;
  LPM_q_ivl_17099 <= tmp_ivl_17101 & tmp_ivl_17096;
  tmp_ivl_17103 <= new_AGEMA_signal_3949 & n3878;
  LPM_q_ivl_17106 <= tmp_ivl_17108 & tmp_ivl_17103;
  new_AGEMA_signal_4276 <= tmp_ivl_17110(1);
  n3518 <= tmp_ivl_17110(0);
  tmp_ivl_17110 <= LPM_d0_ivl_17114(0 + 1 downto 0);
  tmp_ivl_17116 <= z1(54);
  tmp_ivl_17117 <= new_AGEMA_signal_3035 & tmp_ivl_17116;
  LPM_q_ivl_17120 <= tmp_ivl_17122 & tmp_ivl_17117;
  tmp_ivl_17125 <= state_in_s1(270);
  tmp_ivl_17127 <= state_in_s0(270);
  tmp_ivl_17128 <= tmp_ivl_17125 & tmp_ivl_17127;
  LPM_q_ivl_17131 <= tmp_ivl_17133 & tmp_ivl_17128;
  new_AGEMA_signal_3418 <= tmp_ivl_17135(1);
  n3517 <= tmp_ivl_17135(0);
  tmp_ivl_17135 <= LPM_d0_ivl_17139(0 + 1 downto 0);
  tmp_ivl_17141 <= z0(54);
  tmp_ivl_17142 <= new_AGEMA_signal_3226 & tmp_ivl_17141;
  LPM_q_ivl_17145 <= tmp_ivl_17147 & tmp_ivl_17142;
  tmp_ivl_17150 <= state_in_s1(14);
  tmp_ivl_17152 <= state_in_s0(14);
  tmp_ivl_17153 <= tmp_ivl_17150 & tmp_ivl_17152;
  LPM_q_ivl_17156 <= tmp_ivl_17158 & tmp_ivl_17153;
  new_AGEMA_signal_3419 <= tmp_ivl_17160(1);
  n3583 <= tmp_ivl_17160(0);
  tmp_ivl_17160 <= LPM_d0_ivl_17164(0 + 1 downto 0);
  tmp_ivl_17166 <= state_in_s1(78);
  tmp_ivl_17168 <= state_in_s0(78);
  tmp_ivl_17169 <= tmp_ivl_17166 & tmp_ivl_17168;
  LPM_q_ivl_17172 <= tmp_ivl_17174 & tmp_ivl_17169;
  tmp_ivl_17176 <= new_AGEMA_signal_3419 & n3583;
  LPM_q_ivl_17179 <= tmp_ivl_17181 & tmp_ivl_17176;
  new_AGEMA_signal_3701 <= tmp_ivl_17183(1);
  n3516 <= tmp_ivl_17183(0);
  tmp_ivl_17183 <= LPM_d0_ivl_17187(0 + 1 downto 0);
  tmp_ivl_17188 <= new_AGEMA_signal_3418 & n3517;
  LPM_q_ivl_17191 <= tmp_ivl_17193 & tmp_ivl_17188;
  tmp_ivl_17195 <= new_AGEMA_signal_3701 & n3516;
  LPM_q_ivl_17198 <= tmp_ivl_17200 & tmp_ivl_17195;
  new_AGEMA_signal_3978 <= tmp_ivl_17202(1);
  n3524 <= tmp_ivl_17202(0);
  tmp_ivl_17202 <= LPM_d0_ivl_17206(0 + 1 downto 0);
  tmp_ivl_17207 <= new_AGEMA_signal_4276 & n3518;
  LPM_q_ivl_17210 <= tmp_ivl_17212 & tmp_ivl_17207;
  tmp_ivl_17214 <= new_AGEMA_signal_3978 & n3524;
  LPM_q_ivl_17217 <= tmp_ivl_17219 & tmp_ivl_17214;
  tmp_ivl_17221 <= tmp_ivl_17225(1);
  tmp_ivl_17223 <= tmp_ivl_17225(0);
  tmp_ivl_17225 <= LPM_d0_ivl_17229(0 + 1 downto 0);
  tmp_ivl_17230 <= new_AGEMA_signal_3944 & n3519;
  LPM_q_ivl_17233 <= tmp_ivl_17235 & tmp_ivl_17230;
  tmp_ivl_17237 <= new_AGEMA_signal_3978 & n3524;
  LPM_q_ivl_17240 <= tmp_ivl_17242 & tmp_ivl_17237;
  new_AGEMA_signal_4277 <= tmp_ivl_17244(1);
  n3522 <= tmp_ivl_17244(0);
  tmp_ivl_17244 <= LPM_d0_ivl_17248(0 + 1 downto 0);
  tmp_ivl_17250 <= z0(29);
  tmp_ivl_17251 <= new_AGEMA_signal_3259 & tmp_ivl_17250;
  LPM_q_ivl_17254 <= tmp_ivl_17256 & tmp_ivl_17251;
  tmp_ivl_17259 <= state_in_s1(37);
  tmp_ivl_17261 <= state_in_s0(37);
  tmp_ivl_17262 <= tmp_ivl_17259 & tmp_ivl_17261;
  LPM_q_ivl_17265 <= tmp_ivl_17267 & tmp_ivl_17262;
  new_AGEMA_signal_3420 <= tmp_ivl_17269(1);
  n3535 <= tmp_ivl_17269(0);
  tmp_ivl_17269 <= LPM_d0_ivl_17273(0 + 1 downto 0);
  tmp_ivl_17275 <= z1(29);
  tmp_ivl_17276 <= new_AGEMA_signal_3010 & tmp_ivl_17275;
  LPM_q_ivl_17279 <= tmp_ivl_17281 & tmp_ivl_17276;
  tmp_ivl_17283 <= new_AGEMA_signal_3420 & n3535;
  LPM_q_ivl_17286 <= tmp_ivl_17288 & tmp_ivl_17283;
  new_AGEMA_signal_3702 <= tmp_ivl_17290(1);
  n3521 <= tmp_ivl_17290(0);
  tmp_ivl_17290 <= LPM_d0_ivl_17294(0 + 1 downto 0);
  tmp_ivl_17295 <= new_AGEMA_signal_3702 & n3521;
  LPM_q_ivl_17298 <= tmp_ivl_17300 & tmp_ivl_17295;
  tmp_ivl_17302 <= new_AGEMA_signal_2681 & n3520;
  LPM_q_ivl_17305 <= tmp_ivl_17307 & tmp_ivl_17302;
  new_AGEMA_signal_3979 <= tmp_ivl_17309(1);
  n3897 <= tmp_ivl_17309(0);
  tmp_ivl_17309 <= LPM_d0_ivl_17313(0 + 1 downto 0);
  tmp_ivl_17314 <= new_AGEMA_signal_4277 & n3522;
  LPM_q_ivl_17317 <= tmp_ivl_17319 & tmp_ivl_17314;
  tmp_ivl_17321 <= new_AGEMA_signal_3979 & n3897;
  LPM_q_ivl_17324 <= tmp_ivl_17326 & tmp_ivl_17321;
  tmp_ivl_17328 <= tmp_ivl_17332(1);
  tmp_ivl_17330 <= tmp_ivl_17332(0);
  tmp_ivl_17332 <= LPM_d0_ivl_17336(0 + 1 downto 0);
  tmp_ivl_17337 <= new_AGEMA_signal_3971 & n3554;
  LPM_q_ivl_17340 <= tmp_ivl_17342 & tmp_ivl_17337;
  tmp_ivl_17344 <= new_AGEMA_signal_3974 & n3523;
  LPM_q_ivl_17347 <= tmp_ivl_17349 & tmp_ivl_17344;
  new_AGEMA_signal_4278 <= tmp_ivl_17351(1);
  n3525 <= tmp_ivl_17351(0);
  tmp_ivl_17351 <= LPM_d0_ivl_17355(0 + 1 downto 0);
  tmp_ivl_17356 <= new_AGEMA_signal_4278 & n3525;
  LPM_q_ivl_17359 <= tmp_ivl_17361 & tmp_ivl_17356;
  tmp_ivl_17363 <= new_AGEMA_signal_3978 & n3524;
  LPM_q_ivl_17366 <= tmp_ivl_17368 & tmp_ivl_17363;
  tmp_ivl_17370 <= tmp_ivl_17374(1);
  tmp_ivl_17372 <= tmp_ivl_17374(0);
  tmp_ivl_17374 <= LPM_d0_ivl_17378(0 + 1 downto 0);
  tmp_ivl_17380 <= z0(39);
  tmp_ivl_17381 <= new_AGEMA_signal_3222 & tmp_ivl_17380;
  LPM_q_ivl_17384 <= tmp_ivl_17386 & tmp_ivl_17381;
  tmp_ivl_17389 <= state_in_s1(31);
  tmp_ivl_17391 <= state_in_s0(31);
  tmp_ivl_17392 <= tmp_ivl_17389 & tmp_ivl_17391;
  LPM_q_ivl_17395 <= tmp_ivl_17397 & tmp_ivl_17392;
  new_AGEMA_signal_3421 <= tmp_ivl_17399(1);
  n3531 <= tmp_ivl_17399(0);
  tmp_ivl_17399 <= LPM_d0_ivl_17403(0 + 1 downto 0);
  tmp_ivl_17404 <= new_AGEMA_signal_3421 & n3531;
  LPM_q_ivl_17407 <= tmp_ivl_17409 & tmp_ivl_17404;
  tmp_ivl_17411 <= new_AGEMA_signal_3320 & n3526;
  LPM_q_ivl_17414 <= tmp_ivl_17416 & tmp_ivl_17411;
  new_AGEMA_signal_3703 <= tmp_ivl_17418(1);
  n3802 <= tmp_ivl_17418(0);
  tmp_ivl_17418 <= LPM_d0_ivl_17422(0 + 1 downto 0);
  tmp_ivl_17423 <= new_AGEMA_signal_3679 & n3671;
  LPM_q_ivl_17426 <= tmp_ivl_17428 & tmp_ivl_17423;
  tmp_ivl_17430 <= new_AGEMA_signal_3703 & n3802;
  LPM_q_ivl_17433 <= tmp_ivl_17435 & tmp_ivl_17430;
  new_AGEMA_signal_3980 <= tmp_ivl_17437(1);
  n3529 <= tmp_ivl_17437(0);
  tmp_ivl_17437 <= LPM_d0_ivl_17441(0 + 1 downto 0);
  tmp_ivl_17442 <= new_AGEMA_signal_3383 & n3528;
  LPM_q_ivl_17445 <= tmp_ivl_17447 & tmp_ivl_17442;
  tmp_ivl_17449 <= new_AGEMA_signal_3366 & n3527;
  LPM_q_ivl_17452 <= tmp_ivl_17454 & tmp_ivl_17449;
  new_AGEMA_signal_3704 <= tmp_ivl_17456(1);
  n3798 <= tmp_ivl_17456(0);
  tmp_ivl_17456 <= LPM_d0_ivl_17460(0 + 1 downto 0);
  tmp_ivl_17461 <= new_AGEMA_signal_3980 & n3529;
  LPM_q_ivl_17464 <= tmp_ivl_17466 & tmp_ivl_17461;
  tmp_ivl_17468 <= new_AGEMA_signal_3704 & n3798;
  LPM_q_ivl_17471 <= tmp_ivl_17473 & tmp_ivl_17468;
  tmp_ivl_17475 <= tmp_ivl_17479(1);
  tmp_ivl_17477 <= tmp_ivl_17479(0);
  tmp_ivl_17479 <= LPM_d0_ivl_17483(0 + 1 downto 0);
  tmp_ivl_17484 <= new_AGEMA_signal_3959 & n3541;
  LPM_q_ivl_17487 <= tmp_ivl_17489 & tmp_ivl_17484;
  tmp_ivl_17491 <= new_AGEMA_signal_3964 & n3530;
  LPM_q_ivl_17494 <= tmp_ivl_17496 & tmp_ivl_17491;
  new_AGEMA_signal_4280 <= tmp_ivl_17498(1);
  n3534 <= tmp_ivl_17498(0);
  tmp_ivl_17498 <= LPM_d0_ivl_17502(0 + 1 downto 0);
  tmp_ivl_17504 <= z1(39);
  tmp_ivl_17505 <= new_AGEMA_signal_3020 & tmp_ivl_17504;
  LPM_q_ivl_17508 <= tmp_ivl_17510 & tmp_ivl_17505;
  tmp_ivl_17513 <= state_in_s1(287);
  tmp_ivl_17515 <= state_in_s0(287);
  tmp_ivl_17516 <= tmp_ivl_17513 & tmp_ivl_17515;
  LPM_q_ivl_17519 <= tmp_ivl_17521 & tmp_ivl_17516;
  new_AGEMA_signal_3422 <= tmp_ivl_17523(1);
  n3533 <= tmp_ivl_17523(0);
  tmp_ivl_17523 <= LPM_d0_ivl_17527(0 + 1 downto 0);
  tmp_ivl_17529 <= state_in_s1(95);
  tmp_ivl_17531 <= state_in_s0(95);
  tmp_ivl_17532 <= tmp_ivl_17529 & tmp_ivl_17531;
  LPM_q_ivl_17535 <= tmp_ivl_17537 & tmp_ivl_17532;
  tmp_ivl_17539 <= new_AGEMA_signal_3421 & n3531;
  LPM_q_ivl_17542 <= tmp_ivl_17544 & tmp_ivl_17539;
  new_AGEMA_signal_3705 <= tmp_ivl_17546(1);
  n3532 <= tmp_ivl_17546(0);
  tmp_ivl_17546 <= LPM_d0_ivl_17550(0 + 1 downto 0);
  tmp_ivl_17551 <= new_AGEMA_signal_3422 & n3533;
  LPM_q_ivl_17554 <= tmp_ivl_17556 & tmp_ivl_17551;
  tmp_ivl_17558 <= new_AGEMA_signal_3705 & n3532;
  LPM_q_ivl_17561 <= tmp_ivl_17563 & tmp_ivl_17558;
  new_AGEMA_signal_3981 <= tmp_ivl_17565(1);
  n3644 <= tmp_ivl_17565(0);
  tmp_ivl_17565 <= LPM_d0_ivl_17569(0 + 1 downto 0);
  tmp_ivl_17570 <= new_AGEMA_signal_4280 & n3534;
  LPM_q_ivl_17573 <= tmp_ivl_17575 & tmp_ivl_17570;
  tmp_ivl_17577 <= new_AGEMA_signal_3981 & n3644;
  LPM_q_ivl_17580 <= tmp_ivl_17582 & tmp_ivl_17577;
  tmp_ivl_17584 <= tmp_ivl_17588(1);
  tmp_ivl_17586 <= tmp_ivl_17588(0);
  tmp_ivl_17588 <= LPM_d0_ivl_17592(0 + 1 downto 0);
  tmp_ivl_17593 <= new_AGEMA_signal_3697 & n3708;
  LPM_q_ivl_17596 <= tmp_ivl_17598 & tmp_ivl_17593;
  tmp_ivl_17600 <= new_AGEMA_signal_3704 & n3798;
  LPM_q_ivl_17603 <= tmp_ivl_17605 & tmp_ivl_17600;
  new_AGEMA_signal_3982 <= tmp_ivl_17607(1);
  n3536 <= tmp_ivl_17607(0);
  tmp_ivl_17607 <= LPM_d0_ivl_17611(0 + 1 downto 0);
  tmp_ivl_17613 <= state_in_s1(229);
  tmp_ivl_17615 <= state_in_s0(229);
  tmp_ivl_17616 <= tmp_ivl_17613 & tmp_ivl_17615;
  LPM_q_ivl_17619 <= tmp_ivl_17621 & tmp_ivl_17616;
  tmp_ivl_17624 <= z4(29);
  tmp_ivl_17625 <= new_AGEMA_signal_3132 & tmp_ivl_17624;
  LPM_q_ivl_17628 <= tmp_ivl_17630 & tmp_ivl_17625;
  new_AGEMA_signal_3423 <= tmp_ivl_17632(1);
  n3539 <= tmp_ivl_17632(0);
  tmp_ivl_17632 <= LPM_d0_ivl_17636(0 + 1 downto 0);
  tmp_ivl_17637 <= new_AGEMA_signal_3420 & n3535;
  LPM_q_ivl_17640 <= tmp_ivl_17642 & tmp_ivl_17637;
  tmp_ivl_17644 <= new_AGEMA_signal_3423 & n3539;
  LPM_q_ivl_17647 <= tmp_ivl_17649 & tmp_ivl_17644;
  new_AGEMA_signal_3706 <= tmp_ivl_17651(1);
  n3670 <= tmp_ivl_17651(0);
  tmp_ivl_17651 <= LPM_d0_ivl_17655(0 + 1 downto 0);
  tmp_ivl_17656 <= new_AGEMA_signal_3982 & n3536;
  LPM_q_ivl_17659 <= tmp_ivl_17661 & tmp_ivl_17656;
  tmp_ivl_17663 <= new_AGEMA_signal_3706 & n3670;
  LPM_q_ivl_17666 <= tmp_ivl_17668 & tmp_ivl_17663;
  tmp_ivl_17670 <= tmp_ivl_17674(1);
  tmp_ivl_17672 <= tmp_ivl_17674(0);
  tmp_ivl_17674 <= LPM_d0_ivl_17678(0 + 1 downto 0);
  tmp_ivl_17679 <= new_AGEMA_signal_3643 & n3709;
  LPM_q_ivl_17682 <= tmp_ivl_17684 & tmp_ivl_17679;
  tmp_ivl_17686 <= new_AGEMA_signal_3663 & n3843;
  LPM_q_ivl_17689 <= tmp_ivl_17691 & tmp_ivl_17686;
  new_AGEMA_signal_3983 <= tmp_ivl_17693(1);
  n3537 <= tmp_ivl_17693(0);
  tmp_ivl_17693 <= LPM_d0_ivl_17697(0 + 1 downto 0);
  tmp_ivl_17698 <= new_AGEMA_signal_3983 & n3537;
  LPM_q_ivl_17701 <= tmp_ivl_17703 & tmp_ivl_17698;
  tmp_ivl_17705 <= new_AGEMA_signal_3706 & n3670;
  LPM_q_ivl_17708 <= tmp_ivl_17710 & tmp_ivl_17705;
  tmp_ivl_17712 <= tmp_ivl_17716(1);
  tmp_ivl_17714 <= tmp_ivl_17716(0);
  tmp_ivl_17716 <= LPM_d0_ivl_17720(0 + 1 downto 0);
  tmp_ivl_17721 <= new_AGEMA_signal_3609 & n3561;
  LPM_q_ivl_17724 <= tmp_ivl_17726 & tmp_ivl_17721;
  tmp_ivl_17728 <= new_AGEMA_signal_3617 & n3538;
  LPM_q_ivl_17731 <= tmp_ivl_17733 & tmp_ivl_17728;
  new_AGEMA_signal_3984 <= tmp_ivl_17735(1);
  n3540 <= tmp_ivl_17735(0);
  tmp_ivl_17735 <= LPM_d0_ivl_17739(0 + 1 downto 0);
  tmp_ivl_17741 <= state_in_s1(293);
  tmp_ivl_17743 <= state_in_s0(293);
  tmp_ivl_17744 <= tmp_ivl_17741 & tmp_ivl_17743;
  LPM_q_ivl_17747 <= tmp_ivl_17749 & tmp_ivl_17744;
  tmp_ivl_17751 <= new_AGEMA_signal_3423 & n3539;
  LPM_q_ivl_17754 <= tmp_ivl_17756 & tmp_ivl_17751;
  new_AGEMA_signal_3707 <= tmp_ivl_17758(1);
  n3921 <= tmp_ivl_17758(0);
  tmp_ivl_17758 <= LPM_d0_ivl_17762(0 + 1 downto 0);
  tmp_ivl_17763 <= new_AGEMA_signal_3984 & n3540;
  LPM_q_ivl_17766 <= tmp_ivl_17768 & tmp_ivl_17763;
  tmp_ivl_17770 <= new_AGEMA_signal_3707 & n3921;
  LPM_q_ivl_17773 <= tmp_ivl_17775 & tmp_ivl_17770;
  tmp_ivl_17777 <= tmp_ivl_17781(1);
  tmp_ivl_17779 <= tmp_ivl_17781(0);
  tmp_ivl_17781 <= LPM_d0_ivl_17785(0 + 1 downto 0);
  tmp_ivl_17786 <= new_AGEMA_signal_3907 & n3542;
  LPM_q_ivl_17789 <= tmp_ivl_17791 & tmp_ivl_17786;
  tmp_ivl_17793 <= new_AGEMA_signal_3959 & n3541;
  LPM_q_ivl_17796 <= tmp_ivl_17798 & tmp_ivl_17793;
  new_AGEMA_signal_4284 <= tmp_ivl_17800(1);
  n3545 <= tmp_ivl_17800(0);
  tmp_ivl_17800 <= LPM_d0_ivl_17804(0 + 1 downto 0);
  tmp_ivl_17806 <= z1(61);
  tmp_ivl_17807 <= new_AGEMA_signal_3042 & tmp_ivl_17806;
  LPM_q_ivl_17810 <= tmp_ivl_17812 & tmp_ivl_17807;
  tmp_ivl_17815 <= state_in_s1(261);
  tmp_ivl_17817 <= state_in_s0(261);
  tmp_ivl_17818 <= tmp_ivl_17815 & tmp_ivl_17817;
  LPM_q_ivl_17821 <= tmp_ivl_17823 & tmp_ivl_17818;
  new_AGEMA_signal_3424 <= tmp_ivl_17825(1);
  n3544 <= tmp_ivl_17825(0);
  tmp_ivl_17825 <= LPM_d0_ivl_17829(0 + 1 downto 0);
  tmp_ivl_17831 <= z0(61);
  tmp_ivl_17832 <= new_AGEMA_signal_3223 & tmp_ivl_17831;
  LPM_q_ivl_17835 <= tmp_ivl_17837 & tmp_ivl_17832;
  tmp_ivl_17840 <= state_in_s1(5);
  tmp_ivl_17842 <= state_in_s0(5);
  tmp_ivl_17843 <= tmp_ivl_17840 & tmp_ivl_17842;
  LPM_q_ivl_17846 <= tmp_ivl_17848 & tmp_ivl_17843;
  new_AGEMA_signal_3425 <= tmp_ivl_17850(1);
  n3681 <= tmp_ivl_17850(0);
  tmp_ivl_17850 <= LPM_d0_ivl_17854(0 + 1 downto 0);
  tmp_ivl_17856 <= state_in_s1(69);
  tmp_ivl_17858 <= state_in_s0(69);
  tmp_ivl_17859 <= tmp_ivl_17856 & tmp_ivl_17858;
  LPM_q_ivl_17862 <= tmp_ivl_17864 & tmp_ivl_17859;
  tmp_ivl_17866 <= new_AGEMA_signal_3425 & n3681;
  LPM_q_ivl_17869 <= tmp_ivl_17871 & tmp_ivl_17866;
  new_AGEMA_signal_3708 <= tmp_ivl_17873(1);
  n3543 <= tmp_ivl_17873(0);
  tmp_ivl_17873 <= LPM_d0_ivl_17877(0 + 1 downto 0);
  tmp_ivl_17878 <= new_AGEMA_signal_3424 & n3544;
  LPM_q_ivl_17881 <= tmp_ivl_17883 & tmp_ivl_17878;
  tmp_ivl_17885 <= new_AGEMA_signal_3708 & n3543;
  LPM_q_ivl_17888 <= tmp_ivl_17890 & tmp_ivl_17885;
  new_AGEMA_signal_3985 <= tmp_ivl_17892(1);
  n3643 <= tmp_ivl_17892(0);
  tmp_ivl_17892 <= LPM_d0_ivl_17896(0 + 1 downto 0);
  tmp_ivl_17897 <= new_AGEMA_signal_4284 & n3545;
  LPM_q_ivl_17900 <= tmp_ivl_17902 & tmp_ivl_17897;
  tmp_ivl_17904 <= new_AGEMA_signal_3985 & n3643;
  LPM_q_ivl_17907 <= tmp_ivl_17909 & tmp_ivl_17904;
  tmp_ivl_17911 <= tmp_ivl_17915(1);
  tmp_ivl_17913 <= tmp_ivl_17915(0);
  tmp_ivl_17915 <= LPM_d0_ivl_17919(0 + 1 downto 0);
  tmp_ivl_17920 <= new_AGEMA_signal_3921 & n3697;
  LPM_q_ivl_17923 <= tmp_ivl_17925 & tmp_ivl_17920;
  tmp_ivl_17927 <= new_AGEMA_signal_3985 & n3643;
  LPM_q_ivl_17930 <= tmp_ivl_17932 & tmp_ivl_17927;
  new_AGEMA_signal_4285 <= tmp_ivl_17934(1);
  n3549 <= tmp_ivl_17934(0);
  tmp_ivl_17934 <= LPM_d0_ivl_17938(0 + 1 downto 0);
  tmp_ivl_17940 <= z1(22);
  tmp_ivl_17941 <= new_AGEMA_signal_3003 & tmp_ivl_17940;
  LPM_q_ivl_17944 <= tmp_ivl_17946 & tmp_ivl_17941;
  tmp_ivl_17948 <= new_AGEMA_signal_3391 & n3546;
  LPM_q_ivl_17951 <= tmp_ivl_17953 & tmp_ivl_17948;
  new_AGEMA_signal_3709 <= tmp_ivl_17955(1);
  n3548 <= tmp_ivl_17955(0);
  tmp_ivl_17955 <= LPM_d0_ivl_17959(0 + 1 downto 0);
  tmp_ivl_17960 <= new_AGEMA_signal_3709 & n3548;
  LPM_q_ivl_17963 <= tmp_ivl_17965 & tmp_ivl_17960;
  tmp_ivl_17967 <= new_AGEMA_signal_2683 & n3547;
  LPM_q_ivl_17970 <= tmp_ivl_17972 & tmp_ivl_17967;
  new_AGEMA_signal_3986 <= tmp_ivl_17974(1);
  n3702 <= tmp_ivl_17974(0);
  tmp_ivl_17974 <= LPM_d0_ivl_17978(0 + 1 downto 0);
  tmp_ivl_17979 <= new_AGEMA_signal_4285 & n3549;
  LPM_q_ivl_17982 <= tmp_ivl_17984 & tmp_ivl_17979;
  tmp_ivl_17986 <= new_AGEMA_signal_3986 & n3702;
  LPM_q_ivl_17989 <= tmp_ivl_17991 & tmp_ivl_17986;
  tmp_ivl_17993 <= tmp_ivl_17997(1);
  tmp_ivl_17995 <= tmp_ivl_17997(0);
  tmp_ivl_17997 <= LPM_d0_ivl_18001(0 + 1 downto 0);
  tmp_ivl_18003 <= z0(40);
  tmp_ivl_18004 <= new_AGEMA_signal_3220 & tmp_ivl_18003;
  LPM_q_ivl_18007 <= tmp_ivl_18009 & tmp_ivl_18004;
  tmp_ivl_18012 <= state_in_s1(16);
  tmp_ivl_18014 <= state_in_s0(16);
  tmp_ivl_18015 <= tmp_ivl_18012 & tmp_ivl_18014;
  LPM_q_ivl_18018 <= tmp_ivl_18020 & tmp_ivl_18015;
  new_AGEMA_signal_3426 <= tmp_ivl_18022(1);
  n3555 <= tmp_ivl_18022(0);
  tmp_ivl_18022 <= LPM_d0_ivl_18026(0 + 1 downto 0);
  tmp_ivl_18027 <= new_AGEMA_signal_3426 & n3555;
  LPM_q_ivl_18030 <= tmp_ivl_18032 & tmp_ivl_18027;
  tmp_ivl_18034 <= new_AGEMA_signal_3322 & n3550;
  LPM_q_ivl_18037 <= tmp_ivl_18039 & tmp_ivl_18034;
  new_AGEMA_signal_3710 <= tmp_ivl_18041(1);
  n3891 <= tmp_ivl_18041(0);
  tmp_ivl_18041 <= LPM_d0_ivl_18045(0 + 1 downto 0);
  tmp_ivl_18046 <= new_AGEMA_signal_3695 & n3799;
  LPM_q_ivl_18049 <= tmp_ivl_18051 & tmp_ivl_18046;
  tmp_ivl_18053 <= new_AGEMA_signal_3710 & n3891;
  LPM_q_ivl_18056 <= tmp_ivl_18058 & tmp_ivl_18053;
  new_AGEMA_signal_3987 <= tmp_ivl_18060(1);
  n3553 <= tmp_ivl_18060(0);
  tmp_ivl_18060 <= LPM_d0_ivl_18064(0 + 1 downto 0);
  tmp_ivl_18065 <= new_AGEMA_signal_3380 & n3552;
  LPM_q_ivl_18068 <= tmp_ivl_18070 & tmp_ivl_18065;
  tmp_ivl_18072 <= new_AGEMA_signal_3343 & n3551;
  LPM_q_ivl_18075 <= tmp_ivl_18077 & tmp_ivl_18072;
  new_AGEMA_signal_3711 <= tmp_ivl_18079(1);
  n3805 <= tmp_ivl_18079(0);
  tmp_ivl_18079 <= LPM_d0_ivl_18083(0 + 1 downto 0);
  tmp_ivl_18084 <= new_AGEMA_signal_3987 & n3553;
  LPM_q_ivl_18087 <= tmp_ivl_18089 & tmp_ivl_18084;
  tmp_ivl_18091 <= new_AGEMA_signal_3711 & n3805;
  LPM_q_ivl_18094 <= tmp_ivl_18096 & tmp_ivl_18091;
  tmp_ivl_18098 <= tmp_ivl_18102(1);
  tmp_ivl_18100 <= tmp_ivl_18102(0);
  tmp_ivl_18102 <= LPM_d0_ivl_18106(0 + 1 downto 0);
  tmp_ivl_18107 <= new_AGEMA_signal_3971 & n3554;
  LPM_q_ivl_18110 <= tmp_ivl_18112 & tmp_ivl_18107;
  tmp_ivl_18114 <= new_AGEMA_signal_3973 & n3571;
  LPM_q_ivl_18117 <= tmp_ivl_18119 & tmp_ivl_18114;
  new_AGEMA_signal_4287 <= tmp_ivl_18121(1);
  n3558 <= tmp_ivl_18121(0);
  tmp_ivl_18121 <= LPM_d0_ivl_18125(0 + 1 downto 0);
  tmp_ivl_18127 <= z1(40);
  tmp_ivl_18128 <= new_AGEMA_signal_3021 & tmp_ivl_18127;
  LPM_q_ivl_18131 <= tmp_ivl_18133 & tmp_ivl_18128;
  tmp_ivl_18136 <= state_in_s1(272);
  tmp_ivl_18138 <= state_in_s0(272);
  tmp_ivl_18139 <= tmp_ivl_18136 & tmp_ivl_18138;
  LPM_q_ivl_18142 <= tmp_ivl_18144 & tmp_ivl_18139;
  new_AGEMA_signal_3427 <= tmp_ivl_18146(1);
  n3557 <= tmp_ivl_18146(0);
  tmp_ivl_18146 <= LPM_d0_ivl_18150(0 + 1 downto 0);
  tmp_ivl_18152 <= state_in_s1(80);
  tmp_ivl_18154 <= state_in_s0(80);
  tmp_ivl_18155 <= tmp_ivl_18152 & tmp_ivl_18154;
  LPM_q_ivl_18158 <= tmp_ivl_18160 & tmp_ivl_18155;
  tmp_ivl_18162 <= new_AGEMA_signal_3426 & n3555;
  LPM_q_ivl_18165 <= tmp_ivl_18167 & tmp_ivl_18162;
  new_AGEMA_signal_3712 <= tmp_ivl_18169(1);
  n3556 <= tmp_ivl_18169(0);
  tmp_ivl_18169 <= LPM_d0_ivl_18173(0 + 1 downto 0);
  tmp_ivl_18174 <= new_AGEMA_signal_3427 & n3557;
  LPM_q_ivl_18177 <= tmp_ivl_18179 & tmp_ivl_18174;
  tmp_ivl_18181 <= new_AGEMA_signal_3712 & n3556;
  LPM_q_ivl_18184 <= tmp_ivl_18186 & tmp_ivl_18181;
  new_AGEMA_signal_3988 <= tmp_ivl_18188(1);
  n3678 <= tmp_ivl_18188(0);
  tmp_ivl_18188 <= LPM_d0_ivl_18192(0 + 1 downto 0);
  tmp_ivl_18193 <= new_AGEMA_signal_4287 & n3558;
  LPM_q_ivl_18196 <= tmp_ivl_18198 & tmp_ivl_18193;
  tmp_ivl_18200 <= new_AGEMA_signal_3988 & n3678;
  LPM_q_ivl_18203 <= tmp_ivl_18205 & tmp_ivl_18200;
  tmp_ivl_18207 <= tmp_ivl_18211(1);
  tmp_ivl_18209 <= tmp_ivl_18211(0);
  tmp_ivl_18211 <= LPM_d0_ivl_18215(0 + 1 downto 0);
  tmp_ivl_18216 <= new_AGEMA_signal_3587 & n3657;
  LPM_q_ivl_18219 <= tmp_ivl_18221 & tmp_ivl_18216;
  tmp_ivl_18223 <= new_AGEMA_signal_3613 & n3559;
  LPM_q_ivl_18226 <= tmp_ivl_18228 & tmp_ivl_18223;
  new_AGEMA_signal_3989 <= tmp_ivl_18230(1);
  n3560 <= tmp_ivl_18230(0);
  tmp_ivl_18230 <= LPM_d0_ivl_18234(0 + 1 downto 0);
  tmp_ivl_18236 <= state_in_s1(199);
  tmp_ivl_18238 <= state_in_s0(199);
  tmp_ivl_18239 <= tmp_ivl_18236 & tmp_ivl_18238;
  LPM_q_ivl_18242 <= tmp_ivl_18244 & tmp_ivl_18239;
  tmp_ivl_18247 <= z4(63);
  tmp_ivl_18248 <= new_AGEMA_signal_3170 & tmp_ivl_18247;
  LPM_q_ivl_18251 <= tmp_ivl_18253 & tmp_ivl_18248;
  new_AGEMA_signal_3428 <= tmp_ivl_18255(1);
  n3584 <= tmp_ivl_18255(0);
  tmp_ivl_18255 <= LPM_d0_ivl_18259(0 + 1 downto 0);
  tmp_ivl_18261 <= state_in_s1(263);
  tmp_ivl_18263 <= state_in_s0(263);
  tmp_ivl_18264 <= tmp_ivl_18261 & tmp_ivl_18263;
  LPM_q_ivl_18267 <= tmp_ivl_18269 & tmp_ivl_18264;
  tmp_ivl_18271 <= new_AGEMA_signal_3428 & n3584;
  LPM_q_ivl_18274 <= tmp_ivl_18276 & tmp_ivl_18271;
  new_AGEMA_signal_3713 <= tmp_ivl_18278(1);
  n3563 <= tmp_ivl_18278(0);
  tmp_ivl_18278 <= LPM_d0_ivl_18282(0 + 1 downto 0);
  tmp_ivl_18283 <= new_AGEMA_signal_3989 & n3560;
  LPM_q_ivl_18286 <= tmp_ivl_18288 & tmp_ivl_18283;
  tmp_ivl_18290 <= new_AGEMA_signal_3713 & n3563;
  LPM_q_ivl_18293 <= tmp_ivl_18295 & tmp_ivl_18290;
  tmp_ivl_18297 <= tmp_ivl_18301(1);
  tmp_ivl_18299 <= tmp_ivl_18301(0);
  tmp_ivl_18301 <= LPM_d0_ivl_18305(0 + 1 downto 0);
  tmp_ivl_18306 <= new_AGEMA_signal_3609 & n3561;
  LPM_q_ivl_18309 <= tmp_ivl_18311 & tmp_ivl_18306;
  tmp_ivl_18313 <= new_AGEMA_signal_3612 & n3776;
  LPM_q_ivl_18316 <= tmp_ivl_18318 & tmp_ivl_18313;
  new_AGEMA_signal_3990 <= tmp_ivl_18320(1);
  n3562 <= tmp_ivl_18320(0);
  tmp_ivl_18320 <= LPM_d0_ivl_18324(0 + 1 downto 0);
  tmp_ivl_18325 <= new_AGEMA_signal_3990 & n3562;
  LPM_q_ivl_18328 <= tmp_ivl_18330 & tmp_ivl_18325;
  tmp_ivl_18332 <= new_AGEMA_signal_3713 & n3563;
  LPM_q_ivl_18335 <= tmp_ivl_18337 & tmp_ivl_18332;
  tmp_ivl_18339 <= tmp_ivl_18343(1);
  tmp_ivl_18341 <= tmp_ivl_18343(0);
  tmp_ivl_18343 <= LPM_d0_ivl_18347(0 + 1 downto 0);
  tmp_ivl_18348 <= new_AGEMA_signal_3585 & n3926;
  LPM_q_ivl_18351 <= tmp_ivl_18353 & tmp_ivl_18348;
  tmp_ivl_18355 <= new_AGEMA_signal_3707 & n3921;
  LPM_q_ivl_18358 <= tmp_ivl_18360 & tmp_ivl_18355;
  new_AGEMA_signal_3991 <= tmp_ivl_18362(1);
  n3564 <= tmp_ivl_18362(0);
  tmp_ivl_18362 <= LPM_d0_ivl_18366(0 + 1 downto 0);
  tmp_ivl_18367 <= new_AGEMA_signal_3991 & n3564;
  LPM_q_ivl_18370 <= tmp_ivl_18372 & tmp_ivl_18367;
  tmp_ivl_18374 <= new_AGEMA_signal_3713 & n3563;
  LPM_q_ivl_18377 <= tmp_ivl_18379 & tmp_ivl_18374;
  tmp_ivl_18381 <= tmp_ivl_18385(1);
  tmp_ivl_18383 <= tmp_ivl_18385(0);
  tmp_ivl_18385 <= LPM_d0_ivl_18389(0 + 1 downto 0);
  tmp_ivl_18391 <= z0(62);
  tmp_ivl_18392 <= new_AGEMA_signal_3221 & tmp_ivl_18391;
  LPM_q_ivl_18395 <= tmp_ivl_18397 & tmp_ivl_18392;
  tmp_ivl_18400 <= state_in_s1(6);
  tmp_ivl_18402 <= state_in_s0(6);
  tmp_ivl_18403 <= tmp_ivl_18400 & tmp_ivl_18402;
  LPM_q_ivl_18406 <= tmp_ivl_18408 & tmp_ivl_18403;
  new_AGEMA_signal_3429 <= tmp_ivl_18410(1);
  n3573 <= tmp_ivl_18410(0);
  tmp_ivl_18410 <= LPM_d0_ivl_18414(0 + 1 downto 0);
  tmp_ivl_18415 <= new_AGEMA_signal_3429 & n3573;
  LPM_q_ivl_18418 <= tmp_ivl_18420 & tmp_ivl_18415;
  tmp_ivl_18422 <= new_AGEMA_signal_3417 & n3565;
  LPM_q_ivl_18425 <= tmp_ivl_18427 & tmp_ivl_18422;
  new_AGEMA_signal_3714 <= tmp_ivl_18429(1);
  n3872 <= tmp_ivl_18429(0);
  tmp_ivl_18429 <= LPM_d0_ivl_18433(0 + 1 downto 0);
  tmp_ivl_18434 <= new_AGEMA_signal_3407 & n3567;
  LPM_q_ivl_18437 <= tmp_ivl_18439 & tmp_ivl_18434;
  tmp_ivl_18441 <= new_AGEMA_signal_3311 & n3566;
  LPM_q_ivl_18444 <= tmp_ivl_18446 & tmp_ivl_18441;
  new_AGEMA_signal_3715 <= tmp_ivl_18448(1);
  n3773 <= tmp_ivl_18448(0);
  tmp_ivl_18448 <= LPM_d0_ivl_18452(0 + 1 downto 0);
  tmp_ivl_18453 <= new_AGEMA_signal_3714 & n3872;
  LPM_q_ivl_18456 <= tmp_ivl_18458 & tmp_ivl_18453;
  tmp_ivl_18460 <= new_AGEMA_signal_3715 & n3773;
  LPM_q_ivl_18463 <= tmp_ivl_18465 & tmp_ivl_18460;
  new_AGEMA_signal_3992 <= tmp_ivl_18467(1);
  n3570 <= tmp_ivl_18467(0);
  tmp_ivl_18467 <= LPM_d0_ivl_18471(0 + 1 downto 0);
  tmp_ivl_18472 <= new_AGEMA_signal_3339 & n3569;
  LPM_q_ivl_18475 <= tmp_ivl_18477 & tmp_ivl_18472;
  tmp_ivl_18479 <= new_AGEMA_signal_3325 & n3568;
  LPM_q_ivl_18482 <= tmp_ivl_18484 & tmp_ivl_18479;
  new_AGEMA_signal_3716 <= tmp_ivl_18486(1);
  n3760 <= tmp_ivl_18486(0);
  tmp_ivl_18486 <= LPM_d0_ivl_18490(0 + 1 downto 0);
  tmp_ivl_18491 <= new_AGEMA_signal_3992 & n3570;
  LPM_q_ivl_18494 <= tmp_ivl_18496 & tmp_ivl_18491;
  tmp_ivl_18498 <= new_AGEMA_signal_3716 & n3760;
  LPM_q_ivl_18501 <= tmp_ivl_18503 & tmp_ivl_18498;
  tmp_ivl_18505 <= tmp_ivl_18509(1);
  tmp_ivl_18507 <= tmp_ivl_18509(0);
  tmp_ivl_18509 <= LPM_d0_ivl_18513(0 + 1 downto 0);
  tmp_ivl_18514 <= new_AGEMA_signal_3910 & n3572;
  LPM_q_ivl_18517 <= tmp_ivl_18519 & tmp_ivl_18514;
  tmp_ivl_18521 <= new_AGEMA_signal_3973 & n3571;
  LPM_q_ivl_18524 <= tmp_ivl_18526 & tmp_ivl_18521;
  new_AGEMA_signal_4292 <= tmp_ivl_18528(1);
  n3576 <= tmp_ivl_18528(0);
  tmp_ivl_18528 <= LPM_d0_ivl_18532(0 + 1 downto 0);
  tmp_ivl_18534 <= z1(62);
  tmp_ivl_18535 <= new_AGEMA_signal_3043 & tmp_ivl_18534;
  LPM_q_ivl_18538 <= tmp_ivl_18540 & tmp_ivl_18535;
  tmp_ivl_18543 <= state_in_s1(262);
  tmp_ivl_18545 <= state_in_s0(262);
  tmp_ivl_18546 <= tmp_ivl_18543 & tmp_ivl_18545;
  LPM_q_ivl_18549 <= tmp_ivl_18551 & tmp_ivl_18546;
  new_AGEMA_signal_3430 <= tmp_ivl_18553(1);
  n3575 <= tmp_ivl_18553(0);
  tmp_ivl_18553 <= LPM_d0_ivl_18557(0 + 1 downto 0);
  tmp_ivl_18559 <= state_in_s1(70);
  tmp_ivl_18561 <= state_in_s0(70);
  tmp_ivl_18562 <= tmp_ivl_18559 & tmp_ivl_18561;
  LPM_q_ivl_18565 <= tmp_ivl_18567 & tmp_ivl_18562;
  tmp_ivl_18569 <= new_AGEMA_signal_3429 & n3573;
  LPM_q_ivl_18572 <= tmp_ivl_18574 & tmp_ivl_18569;
  new_AGEMA_signal_3717 <= tmp_ivl_18576(1);
  n3574 <= tmp_ivl_18576(0);
  tmp_ivl_18576 <= LPM_d0_ivl_18580(0 + 1 downto 0);
  tmp_ivl_18581 <= new_AGEMA_signal_3430 & n3575;
  LPM_q_ivl_18584 <= tmp_ivl_18586 & tmp_ivl_18581;
  tmp_ivl_18588 <= new_AGEMA_signal_3717 & n3574;
  LPM_q_ivl_18591 <= tmp_ivl_18593 & tmp_ivl_18588;
  new_AGEMA_signal_3993 <= tmp_ivl_18595(1);
  n3677 <= tmp_ivl_18595(0);
  tmp_ivl_18595 <= LPM_d0_ivl_18599(0 + 1 downto 0);
  tmp_ivl_18600 <= new_AGEMA_signal_4292 & n3576;
  LPM_q_ivl_18603 <= tmp_ivl_18605 & tmp_ivl_18600;
  tmp_ivl_18607 <= new_AGEMA_signal_3993 & n3677;
  LPM_q_ivl_18610 <= tmp_ivl_18612 & tmp_ivl_18607;
  tmp_ivl_18614 <= tmp_ivl_18618(1);
  tmp_ivl_18616 <= tmp_ivl_18618(0);
  tmp_ivl_18618 <= LPM_d0_ivl_18622(0 + 1 downto 0);
  tmp_ivl_18623 <= new_AGEMA_signal_3925 & n3796;
  LPM_q_ivl_18626 <= tmp_ivl_18628 & tmp_ivl_18623;
  tmp_ivl_18630 <= new_AGEMA_signal_3993 & n3677;
  LPM_q_ivl_18633 <= tmp_ivl_18635 & tmp_ivl_18630;
  new_AGEMA_signal_4293 <= tmp_ivl_18637(1);
  n3579 <= tmp_ivl_18637(0);
  tmp_ivl_18637 <= LPM_d0_ivl_18641(0 + 1 downto 0);
  tmp_ivl_18643 <= z1(23);
  tmp_ivl_18644 <= new_AGEMA_signal_3004 & tmp_ivl_18643;
  LPM_q_ivl_18647 <= tmp_ivl_18649 & tmp_ivl_18644;
  tmp_ivl_18652 <= state_in_s1(303);
  tmp_ivl_18654 <= state_in_s0(303);
  tmp_ivl_18655 <= tmp_ivl_18652 & tmp_ivl_18654;
  LPM_q_ivl_18658 <= tmp_ivl_18660 & tmp_ivl_18655;
  new_AGEMA_signal_3431 <= tmp_ivl_18662(1);
  n3578 <= tmp_ivl_18662(0);
  tmp_ivl_18662 <= LPM_d0_ivl_18666(0 + 1 downto 0);
  tmp_ivl_18668 <= z0(23);
  tmp_ivl_18669 <= new_AGEMA_signal_3241 & tmp_ivl_18668;
  LPM_q_ivl_18672 <= tmp_ivl_18674 & tmp_ivl_18669;
  tmp_ivl_18677 <= state_in_s1(47);
  tmp_ivl_18679 <= state_in_s0(47);
  tmp_ivl_18680 <= tmp_ivl_18677 & tmp_ivl_18679;
  LPM_q_ivl_18683 <= tmp_ivl_18685 & tmp_ivl_18680;
  new_AGEMA_signal_3432 <= tmp_ivl_18687(1);
  n3595 <= tmp_ivl_18687(0);
  tmp_ivl_18687 <= LPM_d0_ivl_18691(0 + 1 downto 0);
  tmp_ivl_18693 <= state_in_s1(111);
  tmp_ivl_18695 <= state_in_s0(111);
  tmp_ivl_18696 <= tmp_ivl_18693 & tmp_ivl_18695;
  LPM_q_ivl_18699 <= tmp_ivl_18701 & tmp_ivl_18696;
  tmp_ivl_18703 <= new_AGEMA_signal_3432 & n3595;
  LPM_q_ivl_18706 <= tmp_ivl_18708 & tmp_ivl_18703;
  new_AGEMA_signal_3718 <= tmp_ivl_18710(1);
  n3577 <= tmp_ivl_18710(0);
  tmp_ivl_18710 <= LPM_d0_ivl_18714(0 + 1 downto 0);
  tmp_ivl_18715 <= new_AGEMA_signal_3431 & n3578;
  LPM_q_ivl_18718 <= tmp_ivl_18720 & tmp_ivl_18715;
  tmp_ivl_18722 <= new_AGEMA_signal_3718 & n3577;
  LPM_q_ivl_18725 <= tmp_ivl_18727 & tmp_ivl_18722;
  new_AGEMA_signal_3994 <= tmp_ivl_18729(1);
  n3790 <= tmp_ivl_18729(0);
  tmp_ivl_18729 <= LPM_d0_ivl_18733(0 + 1 downto 0);
  tmp_ivl_18734 <= new_AGEMA_signal_4293 & n3579;
  LPM_q_ivl_18737 <= tmp_ivl_18739 & tmp_ivl_18734;
  tmp_ivl_18741 <= new_AGEMA_signal_3994 & n3790;
  LPM_q_ivl_18744 <= tmp_ivl_18746 & tmp_ivl_18741;
  tmp_ivl_18748 <= tmp_ivl_18752(1);
  tmp_ivl_18750 <= tmp_ivl_18752(0);
  tmp_ivl_18752 <= LPM_d0_ivl_18756(0 + 1 downto 0);
  tmp_ivl_18757 <= new_AGEMA_signal_3350 & n3581;
  LPM_q_ivl_18760 <= tmp_ivl_18762 & tmp_ivl_18757;
  tmp_ivl_18764 <= new_AGEMA_signal_3326 & n3580;
  LPM_q_ivl_18767 <= tmp_ivl_18769 & tmp_ivl_18764;
  new_AGEMA_signal_3719 <= tmp_ivl_18771(1);
  n3876 <= tmp_ivl_18771(0);
  tmp_ivl_18771 <= LPM_d0_ivl_18775(0 + 1 downto 0);
  tmp_ivl_18776 <= new_AGEMA_signal_3419 & n3583;
  LPM_q_ivl_18779 <= tmp_ivl_18781 & tmp_ivl_18776;
  tmp_ivl_18783 <= new_AGEMA_signal_3316 & n3582;
  LPM_q_ivl_18786 <= tmp_ivl_18788 & tmp_ivl_18783;
  new_AGEMA_signal_3720 <= tmp_ivl_18790(1);
  n3859 <= tmp_ivl_18790(0);
  tmp_ivl_18790 <= LPM_d0_ivl_18794(0 + 1 downto 0);
  tmp_ivl_18795 <= new_AGEMA_signal_3719 & n3876;
  LPM_q_ivl_18798 <= tmp_ivl_18800 & tmp_ivl_18795;
  tmp_ivl_18802 <= new_AGEMA_signal_3720 & n3859;
  LPM_q_ivl_18805 <= tmp_ivl_18807 & tmp_ivl_18802;
  new_AGEMA_signal_3995 <= tmp_ivl_18809(1);
  n3585 <= tmp_ivl_18809(0);
  tmp_ivl_18809 <= LPM_d0_ivl_18813(0 + 1 downto 0);
  tmp_ivl_18815 <= z0(63);
  tmp_ivl_18816 <= new_AGEMA_signal_3218 & tmp_ivl_18815;
  LPM_q_ivl_18819 <= tmp_ivl_18821 & tmp_ivl_18816;
  tmp_ivl_18824 <= state_in_s1(7);
  tmp_ivl_18826 <= state_in_s0(7);
  tmp_ivl_18827 <= tmp_ivl_18824 & tmp_ivl_18826;
  LPM_q_ivl_18830 <= tmp_ivl_18832 & tmp_ivl_18827;
  new_AGEMA_signal_3433 <= tmp_ivl_18834(1);
  n3587 <= tmp_ivl_18834(0);
  tmp_ivl_18834 <= LPM_d0_ivl_18838(0 + 1 downto 0);
  tmp_ivl_18839 <= new_AGEMA_signal_3433 & n3587;
  LPM_q_ivl_18842 <= tmp_ivl_18844 & tmp_ivl_18839;
  tmp_ivl_18846 <= new_AGEMA_signal_3428 & n3584;
  LPM_q_ivl_18849 <= tmp_ivl_18851 & tmp_ivl_18846;
  new_AGEMA_signal_3721 <= tmp_ivl_18853(1);
  n3855 <= tmp_ivl_18853(0);
  tmp_ivl_18853 <= LPM_d0_ivl_18857(0 + 1 downto 0);
  tmp_ivl_18858 <= new_AGEMA_signal_3995 & n3585;
  LPM_q_ivl_18861 <= tmp_ivl_18863 & tmp_ivl_18858;
  tmp_ivl_18865 <= new_AGEMA_signal_3721 & n3855;
  LPM_q_ivl_18868 <= tmp_ivl_18870 & tmp_ivl_18865;
  tmp_ivl_18872 <= tmp_ivl_18876(1);
  tmp_ivl_18874 <= tmp_ivl_18876(0);
  tmp_ivl_18876 <= LPM_d0_ivl_18880(0 + 1 downto 0);
  tmp_ivl_18881 <= new_AGEMA_signal_3916 & n3586;
  LPM_q_ivl_18884 <= tmp_ivl_18886 & tmp_ivl_18881;
  tmp_ivl_18888 <= new_AGEMA_signal_3951 & n3607;
  LPM_q_ivl_18891 <= tmp_ivl_18893 & tmp_ivl_18888;
  new_AGEMA_signal_4295 <= tmp_ivl_18895(1);
  n3590 <= tmp_ivl_18895(0);
  tmp_ivl_18895 <= LPM_d0_ivl_18899(0 + 1 downto 0);
  tmp_ivl_18901 <= z1(63);
  tmp_ivl_18902 <= new_AGEMA_signal_3044 & tmp_ivl_18901;
  LPM_q_ivl_18905 <= tmp_ivl_18907 & tmp_ivl_18902;
  tmp_ivl_18910 <= state_in_s1(263);
  tmp_ivl_18912 <= state_in_s0(263);
  tmp_ivl_18913 <= tmp_ivl_18910 & tmp_ivl_18912;
  LPM_q_ivl_18916 <= tmp_ivl_18918 & tmp_ivl_18913;
  new_AGEMA_signal_3434 <= tmp_ivl_18920(1);
  n3589 <= tmp_ivl_18920(0);
  tmp_ivl_18920 <= LPM_d0_ivl_18924(0 + 1 downto 0);
  tmp_ivl_18926 <= state_in_s1(71);
  tmp_ivl_18928 <= state_in_s0(71);
  tmp_ivl_18929 <= tmp_ivl_18926 & tmp_ivl_18928;
  LPM_q_ivl_18932 <= tmp_ivl_18934 & tmp_ivl_18929;
  tmp_ivl_18936 <= new_AGEMA_signal_3433 & n3587;
  LPM_q_ivl_18939 <= tmp_ivl_18941 & tmp_ivl_18936;
  new_AGEMA_signal_3722 <= tmp_ivl_18943(1);
  n3588 <= tmp_ivl_18943(0);
  tmp_ivl_18943 <= LPM_d0_ivl_18947(0 + 1 downto 0);
  tmp_ivl_18948 <= new_AGEMA_signal_3434 & n3589;
  LPM_q_ivl_18951 <= tmp_ivl_18953 & tmp_ivl_18948;
  tmp_ivl_18955 <= new_AGEMA_signal_3722 & n3588;
  LPM_q_ivl_18958 <= tmp_ivl_18960 & tmp_ivl_18955;
  new_AGEMA_signal_3996 <= tmp_ivl_18962(1);
  n3720 <= tmp_ivl_18962(0);
  tmp_ivl_18962 <= LPM_d0_ivl_18966(0 + 1 downto 0);
  tmp_ivl_18967 <= new_AGEMA_signal_4295 & n3590;
  LPM_q_ivl_18970 <= tmp_ivl_18972 & tmp_ivl_18967;
  tmp_ivl_18974 <= new_AGEMA_signal_3996 & n3720;
  LPM_q_ivl_18977 <= tmp_ivl_18979 & tmp_ivl_18974;
  tmp_ivl_18981 <= tmp_ivl_18985(1);
  tmp_ivl_18983 <= tmp_ivl_18985(0);
  tmp_ivl_18985 <= LPM_d0_ivl_18989(0 + 1 downto 0);
  tmp_ivl_18990 <= new_AGEMA_signal_3919 & n3853;
  LPM_q_ivl_18993 <= tmp_ivl_18995 & tmp_ivl_18990;
  tmp_ivl_18997 <= new_AGEMA_signal_3996 & n3720;
  LPM_q_ivl_19000 <= tmp_ivl_19002 & tmp_ivl_18997;
  new_AGEMA_signal_4296 <= tmp_ivl_19004(1);
  n3594 <= tmp_ivl_19004(0);
  tmp_ivl_19004 <= LPM_d0_ivl_19008(0 + 1 downto 0);
  tmp_ivl_19010 <= z1(24);
  tmp_ivl_19011 <= new_AGEMA_signal_3005 & tmp_ivl_19010;
  LPM_q_ivl_19014 <= tmp_ivl_19016 & tmp_ivl_19011;
  tmp_ivl_19019 <= state_in_s1(288);
  tmp_ivl_19021 <= state_in_s0(288);
  tmp_ivl_19022 <= tmp_ivl_19019 & tmp_ivl_19021;
  LPM_q_ivl_19025 <= tmp_ivl_19027 & tmp_ivl_19022;
  new_AGEMA_signal_3435 <= tmp_ivl_19029(1);
  n3593 <= tmp_ivl_19029(0);
  tmp_ivl_19029 <= LPM_d0_ivl_19033(0 + 1 downto 0);
  tmp_ivl_19035 <= state_in_s1(96);
  tmp_ivl_19037 <= state_in_s0(96);
  tmp_ivl_19038 <= tmp_ivl_19035 & tmp_ivl_19037;
  LPM_q_ivl_19041 <= tmp_ivl_19043 & tmp_ivl_19038;
  tmp_ivl_19045 <= new_AGEMA_signal_3411 & n3591;
  LPM_q_ivl_19048 <= tmp_ivl_19050 & tmp_ivl_19045;
  new_AGEMA_signal_3723 <= tmp_ivl_19052(1);
  n3592 <= tmp_ivl_19052(0);
  tmp_ivl_19052 <= LPM_d0_ivl_19056(0 + 1 downto 0);
  tmp_ivl_19057 <= new_AGEMA_signal_3435 & n3593;
  LPM_q_ivl_19060 <= tmp_ivl_19062 & tmp_ivl_19057;
  tmp_ivl_19064 <= new_AGEMA_signal_3723 & n3592;
  LPM_q_ivl_19067 <= tmp_ivl_19069 & tmp_ivl_19064;
  new_AGEMA_signal_3997 <= tmp_ivl_19071(1);
  n3848 <= tmp_ivl_19071(0);
  tmp_ivl_19071 <= LPM_d0_ivl_19075(0 + 1 downto 0);
  tmp_ivl_19076 <= new_AGEMA_signal_4296 & n3594;
  LPM_q_ivl_19079 <= tmp_ivl_19081 & tmp_ivl_19076;
  tmp_ivl_19083 <= new_AGEMA_signal_3997 & n3848;
  LPM_q_ivl_19086 <= tmp_ivl_19088 & tmp_ivl_19083;
  tmp_ivl_19090 <= tmp_ivl_19094(1);
  tmp_ivl_19092 <= tmp_ivl_19094(0);
  tmp_ivl_19094 <= LPM_d0_ivl_19098(0 + 1 downto 0);
  tmp_ivl_19100 <= state_in_s1(239);
  tmp_ivl_19102 <= state_in_s0(239);
  tmp_ivl_19103 <= tmp_ivl_19100 & tmp_ivl_19102;
  LPM_q_ivl_19106 <= tmp_ivl_19108 & tmp_ivl_19103;
  tmp_ivl_19111 <= z4(23);
  tmp_ivl_19112 <= new_AGEMA_signal_3126 & tmp_ivl_19111;
  LPM_q_ivl_19115 <= tmp_ivl_19117 & tmp_ivl_19112;
  new_AGEMA_signal_3436 <= tmp_ivl_19119(1);
  n3601 <= tmp_ivl_19119(0);
  tmp_ivl_19119 <= LPM_d0_ivl_19123(0 + 1 downto 0);
  tmp_ivl_19124 <= new_AGEMA_signal_3432 & n3595;
  LPM_q_ivl_19127 <= tmp_ivl_19129 & tmp_ivl_19124;
  tmp_ivl_19131 <= new_AGEMA_signal_3436 & n3601;
  LPM_q_ivl_19134 <= tmp_ivl_19136 & tmp_ivl_19131;
  new_AGEMA_signal_3724 <= tmp_ivl_19138(1);
  n3894 <= tmp_ivl_19138(0);
  tmp_ivl_19138 <= LPM_d0_ivl_19142(0 + 1 downto 0);
  tmp_ivl_19143 <= new_AGEMA_signal_3337 & n3597;
  LPM_q_ivl_19146 <= tmp_ivl_19148 & tmp_ivl_19143;
  tmp_ivl_19150 <= new_AGEMA_signal_3367 & n3596;
  LPM_q_ivl_19153 <= tmp_ivl_19155 & tmp_ivl_19150;
  new_AGEMA_signal_3725 <= tmp_ivl_19157(1);
  n3890 <= tmp_ivl_19157(0);
  tmp_ivl_19157 <= LPM_d0_ivl_19161(0 + 1 downto 0);
  tmp_ivl_19162 <= new_AGEMA_signal_3724 & n3894;
  LPM_q_ivl_19165 <= tmp_ivl_19167 & tmp_ivl_19162;
  tmp_ivl_19169 <= new_AGEMA_signal_3725 & n3890;
  LPM_q_ivl_19172 <= tmp_ivl_19174 & tmp_ivl_19169;
  new_AGEMA_signal_3998 <= tmp_ivl_19176(1);
  n3600 <= tmp_ivl_19176(0);
  tmp_ivl_19176 <= LPM_d0_ivl_19180(0 + 1 downto 0);
  tmp_ivl_19181 <= new_AGEMA_signal_3405 & n3599;
  LPM_q_ivl_19184 <= tmp_ivl_19186 & tmp_ivl_19181;
  tmp_ivl_19188 <= new_AGEMA_signal_3329 & n3598;
  LPM_q_ivl_19191 <= tmp_ivl_19193 & tmp_ivl_19188;
  new_AGEMA_signal_3726 <= tmp_ivl_19195(1);
  n3737 <= tmp_ivl_19195(0);
  tmp_ivl_19195 <= LPM_d0_ivl_19199(0 + 1 downto 0);
  tmp_ivl_19200 <= new_AGEMA_signal_3998 & n3600;
  LPM_q_ivl_19203 <= tmp_ivl_19205 & tmp_ivl_19200;
  tmp_ivl_19207 <= new_AGEMA_signal_3726 & n3737;
  LPM_q_ivl_19210 <= tmp_ivl_19212 & tmp_ivl_19207;
  tmp_ivl_19214 <= tmp_ivl_19218(1);
  tmp_ivl_19216 <= tmp_ivl_19218(0);
  tmp_ivl_19218 <= LPM_d0_ivl_19222(0 + 1 downto 0);
  tmp_ivl_19223 <= new_AGEMA_signal_3601 & n3625;
  LPM_q_ivl_19226 <= tmp_ivl_19228 & tmp_ivl_19223;
  tmp_ivl_19230 <= new_AGEMA_signal_3603 & n3687;
  LPM_q_ivl_19233 <= tmp_ivl_19235 & tmp_ivl_19230;
  new_AGEMA_signal_3999 <= tmp_ivl_19237(1);
  n3602 <= tmp_ivl_19237(0);
  tmp_ivl_19237 <= LPM_d0_ivl_19241(0 + 1 downto 0);
  tmp_ivl_19243 <= state_in_s1(303);
  tmp_ivl_19245 <= state_in_s0(303);
  tmp_ivl_19246 <= tmp_ivl_19243 & tmp_ivl_19245;
  LPM_q_ivl_19249 <= tmp_ivl_19251 & tmp_ivl_19246;
  tmp_ivl_19253 <= new_AGEMA_signal_3436 & n3601;
  LPM_q_ivl_19256 <= tmp_ivl_19258 & tmp_ivl_19253;
  new_AGEMA_signal_3727 <= tmp_ivl_19260(1);
  n3690 <= tmp_ivl_19260(0);
  tmp_ivl_19260 <= LPM_d0_ivl_19264(0 + 1 downto 0);
  tmp_ivl_19265 <= new_AGEMA_signal_3999 & n3602;
  LPM_q_ivl_19268 <= tmp_ivl_19270 & tmp_ivl_19265;
  tmp_ivl_19272 <= new_AGEMA_signal_3727 & n3690;
  LPM_q_ivl_19275 <= tmp_ivl_19277 & tmp_ivl_19272;
  tmp_ivl_19279 <= tmp_ivl_19283(1);
  tmp_ivl_19281 <= tmp_ivl_19283(0);
  tmp_ivl_19283 <= LPM_d0_ivl_19287(0 + 1 downto 0);
  tmp_ivl_19288 <= new_AGEMA_signal_3389 & n3604;
  LPM_q_ivl_19291 <= tmp_ivl_19293 & tmp_ivl_19288;
  tmp_ivl_19295 <= new_AGEMA_signal_3321 & n3603;
  LPM_q_ivl_19298 <= tmp_ivl_19300 & tmp_ivl_19295;
  new_AGEMA_signal_3728 <= tmp_ivl_19302(1);
  n3893 <= tmp_ivl_19302(0);
  tmp_ivl_19302 <= LPM_d0_ivl_19306(0 + 1 downto 0);
  tmp_ivl_19307 <= new_AGEMA_signal_3666 & n3887;
  LPM_q_ivl_19310 <= tmp_ivl_19312 & tmp_ivl_19307;
  tmp_ivl_19314 <= new_AGEMA_signal_3728 & n3893;
  LPM_q_ivl_19317 <= tmp_ivl_19319 & tmp_ivl_19314;
  new_AGEMA_signal_4000 <= tmp_ivl_19321(1);
  n3606 <= tmp_ivl_19321(0);
  tmp_ivl_19321 <= LPM_d0_ivl_19325(0 + 1 downto 0);
  tmp_ivl_19327 <= z0(41);
  tmp_ivl_19328 <= new_AGEMA_signal_3219 & tmp_ivl_19327;
  LPM_q_ivl_19331 <= tmp_ivl_19333 & tmp_ivl_19328;
  tmp_ivl_19336 <= state_in_s1(17);
  tmp_ivl_19338 <= state_in_s0(17);
  tmp_ivl_19339 <= tmp_ivl_19336 & tmp_ivl_19338;
  LPM_q_ivl_19342 <= tmp_ivl_19344 & tmp_ivl_19339;
  new_AGEMA_signal_3437 <= tmp_ivl_19346(1);
  n3609 <= tmp_ivl_19346(0);
  tmp_ivl_19346 <= LPM_d0_ivl_19350(0 + 1 downto 0);
  tmp_ivl_19351 <= new_AGEMA_signal_3437 & n3609;
  LPM_q_ivl_19354 <= tmp_ivl_19356 & tmp_ivl_19351;
  tmp_ivl_19358 <= new_AGEMA_signal_3324 & n3605;
  LPM_q_ivl_19361 <= tmp_ivl_19363 & tmp_ivl_19358;
  new_AGEMA_signal_3729 <= tmp_ivl_19365(1);
  n3740 <= tmp_ivl_19365(0);
  tmp_ivl_19365 <= LPM_d0_ivl_19369(0 + 1 downto 0);
  tmp_ivl_19370 <= new_AGEMA_signal_4000 & n3606;
  LPM_q_ivl_19373 <= tmp_ivl_19375 & tmp_ivl_19370;
  tmp_ivl_19377 <= new_AGEMA_signal_3729 & n3740;
  LPM_q_ivl_19380 <= tmp_ivl_19382 & tmp_ivl_19377;
  tmp_ivl_19384 <= tmp_ivl_19388(1);
  tmp_ivl_19386 <= tmp_ivl_19388(0);
  tmp_ivl_19388 <= LPM_d0_ivl_19392(0 + 1 downto 0);
  tmp_ivl_19393 <= new_AGEMA_signal_3922 & n3608;
  LPM_q_ivl_19396 <= tmp_ivl_19398 & tmp_ivl_19393;
  tmp_ivl_19400 <= new_AGEMA_signal_3951 & n3607;
  LPM_q_ivl_19403 <= tmp_ivl_19405 & tmp_ivl_19400;
  new_AGEMA_signal_4300 <= tmp_ivl_19407(1);
  n3612 <= tmp_ivl_19407(0);
  tmp_ivl_19407 <= LPM_d0_ivl_19411(0 + 1 downto 0);
  tmp_ivl_19413 <= z1(41);
  tmp_ivl_19414 <= new_AGEMA_signal_3022 & tmp_ivl_19413;
  LPM_q_ivl_19417 <= tmp_ivl_19419 & tmp_ivl_19414;
  tmp_ivl_19421 <= new_AGEMA_signal_3437 & n3609;
  LPM_q_ivl_19424 <= tmp_ivl_19426 & tmp_ivl_19421;
  new_AGEMA_signal_3730 <= tmp_ivl_19428(1);
  n3611 <= tmp_ivl_19428(0);
  tmp_ivl_19428 <= LPM_d0_ivl_19432(0 + 1 downto 0);
  tmp_ivl_19433 <= new_AGEMA_signal_3730 & n3611;
  LPM_q_ivl_19436 <= tmp_ivl_19438 & tmp_ivl_19433;
  tmp_ivl_19440 <= new_AGEMA_signal_2685 & n3610;
  LPM_q_ivl_19443 <= tmp_ivl_19445 & tmp_ivl_19440;
  new_AGEMA_signal_4001 <= tmp_ivl_19447(1);
  n3719 <= tmp_ivl_19447(0);
  tmp_ivl_19447 <= LPM_d0_ivl_19451(0 + 1 downto 0);
  tmp_ivl_19452 <= new_AGEMA_signal_4300 & n3612;
  LPM_q_ivl_19455 <= tmp_ivl_19457 & tmp_ivl_19452;
  tmp_ivl_19459 <= new_AGEMA_signal_4001 & n3719;
  LPM_q_ivl_19462 <= tmp_ivl_19464 & tmp_ivl_19459;
  tmp_ivl_19466 <= tmp_ivl_19470(1);
  tmp_ivl_19468 <= tmp_ivl_19470(0);
  tmp_ivl_19470 <= LPM_d0_ivl_19474(0 + 1 downto 0);
  tmp_ivl_19475 <= new_AGEMA_signal_3334 & n3614;
  LPM_q_ivl_19478 <= tmp_ivl_19480 & tmp_ivl_19475;
  tmp_ivl_19482 <= new_AGEMA_signal_3323 & n3613;
  LPM_q_ivl_19485 <= tmp_ivl_19487 & tmp_ivl_19482;
  new_AGEMA_signal_3731 <= tmp_ivl_19489(1);
  n3915 <= tmp_ivl_19489(0);
  tmp_ivl_19489 <= LPM_d0_ivl_19493(0 + 1 downto 0);
  tmp_ivl_19494 <= new_AGEMA_signal_3726 & n3737;
  LPM_q_ivl_19497 <= tmp_ivl_19499 & tmp_ivl_19494;
  tmp_ivl_19501 <= new_AGEMA_signal_3731 & n3915;
  LPM_q_ivl_19504 <= tmp_ivl_19506 & tmp_ivl_19501;
  new_AGEMA_signal_4002 <= tmp_ivl_19508(1);
  n3616 <= tmp_ivl_19508(0);
  tmp_ivl_19508 <= LPM_d0_ivl_19512(0 + 1 downto 0);
  tmp_ivl_19514 <= z0(42);
  tmp_ivl_19515 <= new_AGEMA_signal_3217 & tmp_ivl_19514;
  LPM_q_ivl_19518 <= tmp_ivl_19520 & tmp_ivl_19515;
  tmp_ivl_19523 <= state_in_s1(18);
  tmp_ivl_19525 <= state_in_s0(18);
  tmp_ivl_19526 <= tmp_ivl_19523 & tmp_ivl_19525;
  LPM_q_ivl_19529 <= tmp_ivl_19531 & tmp_ivl_19526;
  new_AGEMA_signal_3438 <= tmp_ivl_19533(1);
  n3618 <= tmp_ivl_19533(0);
  tmp_ivl_19533 <= LPM_d0_ivl_19537(0 + 1 downto 0);
  tmp_ivl_19538 <= new_AGEMA_signal_3438 & n3618;
  LPM_q_ivl_19541 <= tmp_ivl_19543 & tmp_ivl_19538;
  tmp_ivl_19545 <= new_AGEMA_signal_3299 & n3615;
  LPM_q_ivl_19548 <= tmp_ivl_19550 & tmp_ivl_19545;
  new_AGEMA_signal_3732 <= tmp_ivl_19552(1);
  n3828 <= tmp_ivl_19552(0);
  tmp_ivl_19552 <= LPM_d0_ivl_19556(0 + 1 downto 0);
  tmp_ivl_19557 <= new_AGEMA_signal_4002 & n3616;
  LPM_q_ivl_19560 <= tmp_ivl_19562 & tmp_ivl_19557;
  tmp_ivl_19564 <= new_AGEMA_signal_3732 & n3828;
  LPM_q_ivl_19567 <= tmp_ivl_19569 & tmp_ivl_19564;
  tmp_ivl_19571 <= tmp_ivl_19575(1);
  tmp_ivl_19573 <= tmp_ivl_19575(0);
  tmp_ivl_19575 <= LPM_d0_ivl_19579(0 + 1 downto 0);
  tmp_ivl_19580 <= new_AGEMA_signal_3926 & n3617;
  LPM_q_ivl_19583 <= tmp_ivl_19585 & tmp_ivl_19580;
  tmp_ivl_19587 <= new_AGEMA_signal_3981 & n3644;
  LPM_q_ivl_19590 <= tmp_ivl_19592 & tmp_ivl_19587;
  new_AGEMA_signal_4302 <= tmp_ivl_19594(1);
  n3621 <= tmp_ivl_19594(0);
  tmp_ivl_19594 <= LPM_d0_ivl_19598(0 + 1 downto 0);
  tmp_ivl_19600 <= z1(42);
  tmp_ivl_19601 <= new_AGEMA_signal_3023 & tmp_ivl_19600;
  LPM_q_ivl_19604 <= tmp_ivl_19606 & tmp_ivl_19601;
  tmp_ivl_19609 <= state_in_s1(274);
  tmp_ivl_19611 <= state_in_s0(274);
  tmp_ivl_19612 <= tmp_ivl_19609 & tmp_ivl_19611;
  LPM_q_ivl_19615 <= tmp_ivl_19617 & tmp_ivl_19612;
  new_AGEMA_signal_3439 <= tmp_ivl_19619(1);
  n3620 <= tmp_ivl_19619(0);
  tmp_ivl_19619 <= LPM_d0_ivl_19623(0 + 1 downto 0);
  tmp_ivl_19625 <= state_in_s1(82);
  tmp_ivl_19627 <= state_in_s0(82);
  tmp_ivl_19628 <= tmp_ivl_19625 & tmp_ivl_19627;
  LPM_q_ivl_19631 <= tmp_ivl_19633 & tmp_ivl_19628;
  tmp_ivl_19635 <= new_AGEMA_signal_3438 & n3618;
  LPM_q_ivl_19638 <= tmp_ivl_19640 & tmp_ivl_19635;
  new_AGEMA_signal_3733 <= tmp_ivl_19642(1);
  n3619 <= tmp_ivl_19642(0);
  tmp_ivl_19642 <= LPM_d0_ivl_19646(0 + 1 downto 0);
  tmp_ivl_19647 <= new_AGEMA_signal_3439 & n3620;
  LPM_q_ivl_19650 <= tmp_ivl_19652 & tmp_ivl_19647;
  tmp_ivl_19654 <= new_AGEMA_signal_3733 & n3619;
  LPM_q_ivl_19657 <= tmp_ivl_19659 & tmp_ivl_19654;
  new_AGEMA_signal_4003 <= tmp_ivl_19661(1);
  n3816 <= tmp_ivl_19661(0);
  tmp_ivl_19661 <= LPM_d0_ivl_19665(0 + 1 downto 0);
  tmp_ivl_19666 <= new_AGEMA_signal_4302 & n3621;
  LPM_q_ivl_19669 <= tmp_ivl_19671 & tmp_ivl_19666;
  tmp_ivl_19673 <= new_AGEMA_signal_4003 & n3816;
  LPM_q_ivl_19676 <= tmp_ivl_19678 & tmp_ivl_19673;
  tmp_ivl_19680 <= tmp_ivl_19684(1);
  tmp_ivl_19682 <= tmp_ivl_19684(0);
  tmp_ivl_19684 <= LPM_d0_ivl_19688(0 + 1 downto 0);
  tmp_ivl_19689 <= new_AGEMA_signal_3678 & n3704;
  LPM_q_ivl_19692 <= tmp_ivl_19694 & tmp_ivl_19689;
  tmp_ivl_19696 <= new_AGEMA_signal_3703 & n3802;
  LPM_q_ivl_19699 <= tmp_ivl_19701 & tmp_ivl_19696;
  new_AGEMA_signal_4004 <= tmp_ivl_19703(1);
  n3623 <= tmp_ivl_19703(0);
  tmp_ivl_19703 <= LPM_d0_ivl_19707(0 + 1 downto 0);
  tmp_ivl_19709 <= state_in_s1(230);
  tmp_ivl_19711 <= state_in_s0(230);
  tmp_ivl_19712 <= tmp_ivl_19709 & tmp_ivl_19711;
  LPM_q_ivl_19715 <= tmp_ivl_19717 & tmp_ivl_19712;
  tmp_ivl_19720 <= z4(30);
  tmp_ivl_19721 <= new_AGEMA_signal_3134 & tmp_ivl_19720;
  LPM_q_ivl_19724 <= tmp_ivl_19726 & tmp_ivl_19721;
  new_AGEMA_signal_3440 <= tmp_ivl_19728(1);
  n3626 <= tmp_ivl_19728(0);
  tmp_ivl_19728 <= LPM_d0_ivl_19732(0 + 1 downto 0);
  tmp_ivl_19733 <= new_AGEMA_signal_3371 & n3622;
  LPM_q_ivl_19736 <= tmp_ivl_19738 & tmp_ivl_19733;
  tmp_ivl_19740 <= new_AGEMA_signal_3440 & n3626;
  LPM_q_ivl_19743 <= tmp_ivl_19745 & tmp_ivl_19740;
  new_AGEMA_signal_3734 <= tmp_ivl_19747(1);
  n3711 <= tmp_ivl_19747(0);
  tmp_ivl_19747 <= LPM_d0_ivl_19751(0 + 1 downto 0);
  tmp_ivl_19752 <= new_AGEMA_signal_4004 & n3623;
  LPM_q_ivl_19755 <= tmp_ivl_19757 & tmp_ivl_19752;
  tmp_ivl_19759 <= new_AGEMA_signal_3734 & n3711;
  LPM_q_ivl_19762 <= tmp_ivl_19764 & tmp_ivl_19759;
  tmp_ivl_19766 <= tmp_ivl_19770(1);
  tmp_ivl_19768 <= tmp_ivl_19770(0);
  tmp_ivl_19770 <= LPM_d0_ivl_19774(0 + 1 downto 0);
  tmp_ivl_19775 <= new_AGEMA_signal_3601 & n3625;
  LPM_q_ivl_19778 <= tmp_ivl_19780 & tmp_ivl_19775;
  tmp_ivl_19782 <= new_AGEMA_signal_3661 & n3624;
  LPM_q_ivl_19785 <= tmp_ivl_19787 & tmp_ivl_19782;
  new_AGEMA_signal_4005 <= tmp_ivl_19789(1);
  n3627 <= tmp_ivl_19789(0);
  tmp_ivl_19789 <= LPM_d0_ivl_19793(0 + 1 downto 0);
  tmp_ivl_19795 <= state_in_s1(294);
  tmp_ivl_19797 <= state_in_s0(294);
  tmp_ivl_19798 <= tmp_ivl_19795 & tmp_ivl_19797;
  LPM_q_ivl_19801 <= tmp_ivl_19803 & tmp_ivl_19798;
  tmp_ivl_19805 <= new_AGEMA_signal_3440 & n3626;
  LPM_q_ivl_19808 <= tmp_ivl_19810 & tmp_ivl_19805;
  new_AGEMA_signal_3735 <= tmp_ivl_19812(1);
  n3632 <= tmp_ivl_19812(0);
  tmp_ivl_19812 <= LPM_d0_ivl_19816(0 + 1 downto 0);
  tmp_ivl_19817 <= new_AGEMA_signal_4005 & n3627;
  LPM_q_ivl_19820 <= tmp_ivl_19822 & tmp_ivl_19817;
  tmp_ivl_19824 <= new_AGEMA_signal_3735 & n3632;
  LPM_q_ivl_19827 <= tmp_ivl_19829 & tmp_ivl_19824;
  tmp_ivl_19831 <= tmp_ivl_19835(1);
  tmp_ivl_19833 <= tmp_ivl_19835(0);
  tmp_ivl_19835 <= LPM_d0_ivl_19839(0 + 1 downto 0);
  tmp_ivl_19840 <= new_AGEMA_signal_3618 & n3629;
  LPM_q_ivl_19843 <= tmp_ivl_19845 & tmp_ivl_19840;
  tmp_ivl_19847 <= new_AGEMA_signal_3655 & n3628;
  LPM_q_ivl_19850 <= tmp_ivl_19852 & tmp_ivl_19847;
  new_AGEMA_signal_4006 <= tmp_ivl_19854(1);
  n3630 <= tmp_ivl_19854(0);
  tmp_ivl_19854 <= LPM_d0_ivl_19858(0 + 1 downto 0);
  tmp_ivl_19859 <= new_AGEMA_signal_4006 & n3630;
  LPM_q_ivl_19862 <= tmp_ivl_19864 & tmp_ivl_19859;
  tmp_ivl_19866 <= new_AGEMA_signal_3735 & n3632;
  LPM_q_ivl_19869 <= tmp_ivl_19871 & tmp_ivl_19866;
  tmp_ivl_19873 <= tmp_ivl_19877(1);
  tmp_ivl_19875 <= tmp_ivl_19877(0);
  tmp_ivl_19877 <= LPM_d0_ivl_19881(0 + 1 downto 0);
  tmp_ivl_19882 <= new_AGEMA_signal_3631 & n3631;
  LPM_q_ivl_19885 <= tmp_ivl_19887 & tmp_ivl_19882;
  tmp_ivl_19889 <= new_AGEMA_signal_3727 & n3690;
  LPM_q_ivl_19892 <= tmp_ivl_19894 & tmp_ivl_19889;
  new_AGEMA_signal_4007 <= tmp_ivl_19896(1);
  n3633 <= tmp_ivl_19896(0);
  tmp_ivl_19896 <= LPM_d0_ivl_19900(0 + 1 downto 0);
  tmp_ivl_19901 <= new_AGEMA_signal_4007 & n3633;
  LPM_q_ivl_19904 <= tmp_ivl_19906 & tmp_ivl_19901;
  tmp_ivl_19908 <= new_AGEMA_signal_3735 & n3632;
  LPM_q_ivl_19911 <= tmp_ivl_19913 & tmp_ivl_19908;
  tmp_ivl_19915 <= tmp_ivl_19919(1);
  tmp_ivl_19917 <= tmp_ivl_19919(0);
  tmp_ivl_19919 <= LPM_d0_ivl_19923(0 + 1 downto 0);
  tmp_ivl_19924 <= new_AGEMA_signal_3662 & n3846;
  LPM_q_ivl_19927 <= tmp_ivl_19929 & tmp_ivl_19924;
  tmp_ivl_19931 <= new_AGEMA_signal_3672 & n3787;
  LPM_q_ivl_19934 <= tmp_ivl_19936 & tmp_ivl_19931;
  new_AGEMA_signal_4008 <= tmp_ivl_19938(1);
  n3635 <= tmp_ivl_19938(0);
  tmp_ivl_19938 <= LPM_d0_ivl_19942(0 + 1 downto 0);
  tmp_ivl_19944 <= z0(0);
  tmp_ivl_19945 <= new_AGEMA_signal_3584 & tmp_ivl_19944;
  LPM_q_ivl_19948 <= tmp_ivl_19950 & tmp_ivl_19945;
  tmp_ivl_19953 <= state_in_s1(56);
  tmp_ivl_19955 <= state_in_s0(56);
  tmp_ivl_19956 <= tmp_ivl_19953 & tmp_ivl_19955;
  LPM_q_ivl_19959 <= tmp_ivl_19961 & tmp_ivl_19956;
  new_AGEMA_signal_3736 <= tmp_ivl_19963(1);
  n3639 <= tmp_ivl_19963(0);
  tmp_ivl_19963 <= LPM_d0_ivl_19967(0 + 1 downto 0);
  tmp_ivl_19968 <= new_AGEMA_signal_3736 & n3639;
  LPM_q_ivl_19971 <= tmp_ivl_19973 & tmp_ivl_19968;
  tmp_ivl_19975 <= new_AGEMA_signal_3345 & n3634;
  LPM_q_ivl_19978 <= tmp_ivl_19980 & tmp_ivl_19975;
  new_AGEMA_signal_4009 <= tmp_ivl_19982(1);
  n3782 <= tmp_ivl_19982(0);
  tmp_ivl_19982 <= LPM_d0_ivl_19986(0 + 1 downto 0);
  tmp_ivl_19987 <= new_AGEMA_signal_4008 & n3635;
  LPM_q_ivl_19990 <= tmp_ivl_19992 & tmp_ivl_19987;
  tmp_ivl_19994 <= new_AGEMA_signal_4009 & n3782;
  LPM_q_ivl_19997 <= tmp_ivl_19999 & tmp_ivl_19994;
  tmp_ivl_20001 <= tmp_ivl_20005(1);
  tmp_ivl_20003 <= tmp_ivl_20005(0);
  tmp_ivl_20005 <= LPM_d0_ivl_20009(0 + 1 downto 0);
  tmp_ivl_20010 <= new_AGEMA_signal_3645 & n3637;
  LPM_q_ivl_20013 <= tmp_ivl_20015 & tmp_ivl_20010;
  tmp_ivl_20017 <= new_AGEMA_signal_3687 & n3636;
  LPM_q_ivl_20020 <= tmp_ivl_20022 & tmp_ivl_20017;
  new_AGEMA_signal_4010 <= tmp_ivl_20024(1);
  n3638 <= tmp_ivl_20024(0);
  tmp_ivl_20024 <= LPM_d0_ivl_20028(0 + 1 downto 0);
  tmp_ivl_20029 <= new_AGEMA_signal_4010 & n3638;
  LPM_q_ivl_20032 <= tmp_ivl_20034 & tmp_ivl_20029;
  tmp_ivl_20036 <= new_AGEMA_signal_4009 & n3782;
  LPM_q_ivl_20039 <= tmp_ivl_20041 & tmp_ivl_20036;
  tmp_ivl_20043 <= tmp_ivl_20047(1);
  tmp_ivl_20045 <= tmp_ivl_20047(0);
  tmp_ivl_20047 <= LPM_d0_ivl_20051(0 + 1 downto 0);
  tmp_ivl_20052 <= new_AGEMA_signal_3934 & n3810;
  LPM_q_ivl_20055 <= tmp_ivl_20057 & tmp_ivl_20052;
  tmp_ivl_20059 <= new_AGEMA_signal_3986 & n3702;
  LPM_q_ivl_20062 <= tmp_ivl_20064 & tmp_ivl_20059;
  new_AGEMA_signal_4309 <= tmp_ivl_20066(1);
  n3642 <= tmp_ivl_20066(0);
  tmp_ivl_20066 <= LPM_d0_ivl_20070(0 + 1 downto 0);
  tmp_ivl_20072 <= z1(0);
  tmp_ivl_20073 <= new_AGEMA_signal_3517 & tmp_ivl_20072;
  LPM_q_ivl_20076 <= tmp_ivl_20078 & tmp_ivl_20073;
  tmp_ivl_20081 <= state_in_s1(312);
  tmp_ivl_20083 <= state_in_s0(312);
  tmp_ivl_20084 <= tmp_ivl_20081 & tmp_ivl_20083;
  LPM_q_ivl_20087 <= tmp_ivl_20089 & tmp_ivl_20084;
  new_AGEMA_signal_3737 <= tmp_ivl_20091(1);
  n3641 <= tmp_ivl_20091(0);
  tmp_ivl_20091 <= LPM_d0_ivl_20095(0 + 1 downto 0);
  tmp_ivl_20097 <= state_in_s1(120);
  tmp_ivl_20099 <= state_in_s0(120);
  tmp_ivl_20100 <= tmp_ivl_20097 & tmp_ivl_20099;
  LPM_q_ivl_20103 <= tmp_ivl_20105 & tmp_ivl_20100;
  tmp_ivl_20107 <= new_AGEMA_signal_3736 & n3639;
  LPM_q_ivl_20110 <= tmp_ivl_20112 & tmp_ivl_20107;
  new_AGEMA_signal_4011 <= tmp_ivl_20114(1);
  n3640 <= tmp_ivl_20114(0);
  tmp_ivl_20114 <= LPM_d0_ivl_20118(0 + 1 downto 0);
  tmp_ivl_20119 <= new_AGEMA_signal_3737 & n3641;
  LPM_q_ivl_20122 <= tmp_ivl_20124 & tmp_ivl_20119;
  tmp_ivl_20126 <= new_AGEMA_signal_4011 & n3640;
  LPM_q_ivl_20129 <= tmp_ivl_20131 & tmp_ivl_20126;
  new_AGEMA_signal_4310 <= tmp_ivl_20133(1);
  n3815 <= tmp_ivl_20133(0);
  tmp_ivl_20133 <= LPM_d0_ivl_20137(0 + 1 downto 0);
  tmp_ivl_20138 <= new_AGEMA_signal_4309 & n3642;
  LPM_q_ivl_20141 <= tmp_ivl_20143 & tmp_ivl_20138;
  tmp_ivl_20145 <= new_AGEMA_signal_4310 & n3815;
  LPM_q_ivl_20148 <= tmp_ivl_20150 & tmp_ivl_20145;
  tmp_ivl_20152 <= tmp_ivl_20156(1);
  tmp_ivl_20154 <= tmp_ivl_20156(0);
  tmp_ivl_20156 <= LPM_d0_ivl_20160(0 + 1 downto 0);
  tmp_ivl_20161 <= new_AGEMA_signal_3981 & n3644;
  LPM_q_ivl_20164 <= tmp_ivl_20166 & tmp_ivl_20161;
  tmp_ivl_20168 <= new_AGEMA_signal_3985 & n3643;
  LPM_q_ivl_20171 <= tmp_ivl_20173 & tmp_ivl_20168;
  new_AGEMA_signal_4311 <= tmp_ivl_20175(1);
  n3645 <= tmp_ivl_20175(0);
  tmp_ivl_20175 <= LPM_d0_ivl_20179(0 + 1 downto 0);
  tmp_ivl_20180 <= new_AGEMA_signal_4311 & n3645;
  LPM_q_ivl_20183 <= tmp_ivl_20185 & tmp_ivl_20180;
  tmp_ivl_20187 <= new_AGEMA_signal_4310 & n3815;
  LPM_q_ivl_20190 <= tmp_ivl_20192 & tmp_ivl_20187;
  tmp_ivl_20194 <= tmp_ivl_20198(1);
  tmp_ivl_20196 <= tmp_ivl_20198(0);
  tmp_ivl_20198 <= LPM_d0_ivl_20202(0 + 1 downto 0);
  tmp_ivl_20203 <= new_AGEMA_signal_3693 & n3823;
  LPM_q_ivl_20206 <= tmp_ivl_20208 & tmp_ivl_20203;
  tmp_ivl_20210 <= new_AGEMA_signal_3716 & n3760;
  LPM_q_ivl_20213 <= tmp_ivl_20215 & tmp_ivl_20210;
  new_AGEMA_signal_4012 <= tmp_ivl_20217(1);
  n3647 <= tmp_ivl_20217(0);
  tmp_ivl_20217 <= LPM_d0_ivl_20221(0 + 1 downto 0);
  tmp_ivl_20223 <= z0(43);
  tmp_ivl_20224 <= new_AGEMA_signal_3216 & tmp_ivl_20223;
  LPM_q_ivl_20227 <= tmp_ivl_20229 & tmp_ivl_20224;
  tmp_ivl_20232 <= state_in_s1(19);
  tmp_ivl_20234 <= state_in_s0(19);
  tmp_ivl_20235 <= tmp_ivl_20232 & tmp_ivl_20234;
  LPM_q_ivl_20238 <= tmp_ivl_20240 & tmp_ivl_20235;
  new_AGEMA_signal_3441 <= tmp_ivl_20242(1);
  n3649 <= tmp_ivl_20242(0);
  tmp_ivl_20242 <= LPM_d0_ivl_20246(0 + 1 downto 0);
  tmp_ivl_20247 <= new_AGEMA_signal_3441 & n3649;
  LPM_q_ivl_20250 <= tmp_ivl_20252 & tmp_ivl_20247;
  tmp_ivl_20254 <= new_AGEMA_signal_3302 & n3646;
  LPM_q_ivl_20257 <= tmp_ivl_20259 & tmp_ivl_20254;
  new_AGEMA_signal_3738 <= tmp_ivl_20261(1);
  n3917 <= tmp_ivl_20261(0);
  tmp_ivl_20261 <= LPM_d0_ivl_20265(0 + 1 downto 0);
  tmp_ivl_20266 <= new_AGEMA_signal_4012 & n3647;
  LPM_q_ivl_20269 <= tmp_ivl_20271 & tmp_ivl_20266;
  tmp_ivl_20273 <= new_AGEMA_signal_3738 & n3917;
  LPM_q_ivl_20276 <= tmp_ivl_20278 & tmp_ivl_20273;
  tmp_ivl_20280 <= tmp_ivl_20284(1);
  tmp_ivl_20282 <= tmp_ivl_20284(0);
  tmp_ivl_20284 <= LPM_d0_ivl_20288(0 + 1 downto 0);
  tmp_ivl_20289 <= new_AGEMA_signal_3920 & n3648;
  LPM_q_ivl_20292 <= tmp_ivl_20294 & tmp_ivl_20289;
  tmp_ivl_20296 <= new_AGEMA_signal_3988 & n3678;
  LPM_q_ivl_20299 <= tmp_ivl_20301 & tmp_ivl_20296;
  new_AGEMA_signal_4313 <= tmp_ivl_20303(1);
  n3652 <= tmp_ivl_20303(0);
  tmp_ivl_20303 <= LPM_d0_ivl_20307(0 + 1 downto 0);
  tmp_ivl_20309 <= z1(43);
  tmp_ivl_20310 <= new_AGEMA_signal_3024 & tmp_ivl_20309;
  LPM_q_ivl_20313 <= tmp_ivl_20315 & tmp_ivl_20310;
  tmp_ivl_20318 <= state_in_s1(275);
  tmp_ivl_20320 <= state_in_s0(275);
  tmp_ivl_20321 <= tmp_ivl_20318 & tmp_ivl_20320;
  LPM_q_ivl_20324 <= tmp_ivl_20326 & tmp_ivl_20321;
  new_AGEMA_signal_3442 <= tmp_ivl_20328(1);
  n3651 <= tmp_ivl_20328(0);
  tmp_ivl_20328 <= LPM_d0_ivl_20332(0 + 1 downto 0);
  tmp_ivl_20334 <= state_in_s1(83);
  tmp_ivl_20336 <= state_in_s0(83);
  tmp_ivl_20337 <= tmp_ivl_20334 & tmp_ivl_20336;
  LPM_q_ivl_20340 <= tmp_ivl_20342 & tmp_ivl_20337;
  tmp_ivl_20344 <= new_AGEMA_signal_3441 & n3649;
  LPM_q_ivl_20347 <= tmp_ivl_20349 & tmp_ivl_20344;
  new_AGEMA_signal_3739 <= tmp_ivl_20351(1);
  n3650 <= tmp_ivl_20351(0);
  tmp_ivl_20351 <= LPM_d0_ivl_20355(0 + 1 downto 0);
  tmp_ivl_20356 <= new_AGEMA_signal_3442 & n3651;
  LPM_q_ivl_20359 <= tmp_ivl_20361 & tmp_ivl_20356;
  tmp_ivl_20363 <= new_AGEMA_signal_3739 & n3650;
  LPM_q_ivl_20366 <= tmp_ivl_20368 & tmp_ivl_20363;
  new_AGEMA_signal_4013 <= tmp_ivl_20370(1);
  n3904 <= tmp_ivl_20370(0);
  tmp_ivl_20370 <= LPM_d0_ivl_20374(0 + 1 downto 0);
  tmp_ivl_20375 <= new_AGEMA_signal_4313 & n3652;
  LPM_q_ivl_20378 <= tmp_ivl_20380 & tmp_ivl_20375;
  tmp_ivl_20382 <= new_AGEMA_signal_4013 & n3904;
  LPM_q_ivl_20385 <= tmp_ivl_20387 & tmp_ivl_20382;
  tmp_ivl_20389 <= tmp_ivl_20393(1);
  tmp_ivl_20391 <= tmp_ivl_20393(0);
  tmp_ivl_20393 <= LPM_d0_ivl_20397(0 + 1 downto 0);
  tmp_ivl_20398 <= new_AGEMA_signal_3668 & n3803;
  LPM_q_ivl_20401 <= tmp_ivl_20403 & tmp_ivl_20398;
  tmp_ivl_20405 <= new_AGEMA_signal_3734 & n3711;
  LPM_q_ivl_20408 <= tmp_ivl_20410 & tmp_ivl_20405;
  new_AGEMA_signal_4014 <= tmp_ivl_20412(1);
  n3654 <= tmp_ivl_20412(0);
  tmp_ivl_20412 <= LPM_d0_ivl_20416(0 + 1 downto 0);
  tmp_ivl_20418 <= state_in_s1(201);
  tmp_ivl_20420 <= state_in_s0(201);
  tmp_ivl_20421 <= tmp_ivl_20418 & tmp_ivl_20420;
  LPM_q_ivl_20424 <= tmp_ivl_20426 & tmp_ivl_20421;
  tmp_ivl_20429 <= z4(49);
  tmp_ivl_20430 <= new_AGEMA_signal_3154 & tmp_ivl_20429;
  LPM_q_ivl_20433 <= tmp_ivl_20435 & tmp_ivl_20430;
  new_AGEMA_signal_3443 <= tmp_ivl_20437(1);
  n3658 <= tmp_ivl_20437(0);
  tmp_ivl_20437 <= LPM_d0_ivl_20441(0 + 1 downto 0);
  tmp_ivl_20442 <= new_AGEMA_signal_3398 & n3653;
  LPM_q_ivl_20445 <= tmp_ivl_20447 & tmp_ivl_20442;
  tmp_ivl_20449 <= new_AGEMA_signal_3443 & n3658;
  LPM_q_ivl_20452 <= tmp_ivl_20454 & tmp_ivl_20449;
  new_AGEMA_signal_3740 <= tmp_ivl_20456(1);
  n3886 <= tmp_ivl_20456(0);
  tmp_ivl_20456 <= LPM_d0_ivl_20460(0 + 1 downto 0);
  tmp_ivl_20461 <= new_AGEMA_signal_4014 & n3654;
  LPM_q_ivl_20464 <= tmp_ivl_20466 & tmp_ivl_20461;
  tmp_ivl_20468 <= new_AGEMA_signal_3740 & n3886;
  LPM_q_ivl_20471 <= tmp_ivl_20473 & tmp_ivl_20468;
  tmp_ivl_20475 <= tmp_ivl_20479(1);
  tmp_ivl_20477 <= tmp_ivl_20479(0);
  tmp_ivl_20479 <= LPM_d0_ivl_20483(0 + 1 downto 0);
  tmp_ivl_20484 <= new_AGEMA_signal_3696 & n3712;
  LPM_q_ivl_20487 <= tmp_ivl_20489 & tmp_ivl_20484;
  tmp_ivl_20491 <= new_AGEMA_signal_3710 & n3891;
  LPM_q_ivl_20494 <= tmp_ivl_20496 & tmp_ivl_20491;
  new_AGEMA_signal_4015 <= tmp_ivl_20498(1);
  n3655 <= tmp_ivl_20498(0);
  tmp_ivl_20498 <= LPM_d0_ivl_20502(0 + 1 downto 0);
  tmp_ivl_20503 <= new_AGEMA_signal_4015 & n3655;
  LPM_q_ivl_20506 <= tmp_ivl_20508 & tmp_ivl_20503;
  tmp_ivl_20510 <= new_AGEMA_signal_3740 & n3886;
  LPM_q_ivl_20513 <= tmp_ivl_20515 & tmp_ivl_20510;
  tmp_ivl_20517 <= tmp_ivl_20521(1);
  tmp_ivl_20519 <= tmp_ivl_20521(0);
  tmp_ivl_20521 <= LPM_d0_ivl_20525(0 + 1 downto 0);
  tmp_ivl_20526 <= new_AGEMA_signal_3587 & n3657;
  LPM_q_ivl_20529 <= tmp_ivl_20531 & tmp_ivl_20526;
  tmp_ivl_20533 <= new_AGEMA_signal_3654 & n3656;
  LPM_q_ivl_20536 <= tmp_ivl_20538 & tmp_ivl_20533;
  new_AGEMA_signal_4016 <= tmp_ivl_20540(1);
  n3659 <= tmp_ivl_20540(0);
  tmp_ivl_20540 <= LPM_d0_ivl_20544(0 + 1 downto 0);
  tmp_ivl_20546 <= state_in_s1(265);
  tmp_ivl_20548 <= state_in_s0(265);
  tmp_ivl_20549 <= tmp_ivl_20546 & tmp_ivl_20548;
  LPM_q_ivl_20552 <= tmp_ivl_20554 & tmp_ivl_20549;
  tmp_ivl_20556 <= new_AGEMA_signal_3443 & n3658;
  LPM_q_ivl_20559 <= tmp_ivl_20561 & tmp_ivl_20556;
  new_AGEMA_signal_3741 <= tmp_ivl_20563(1);
  n3665 <= tmp_ivl_20563(0);
  tmp_ivl_20563 <= LPM_d0_ivl_20567(0 + 1 downto 0);
  tmp_ivl_20568 <= new_AGEMA_signal_4016 & n3659;
  LPM_q_ivl_20571 <= tmp_ivl_20573 & tmp_ivl_20568;
  tmp_ivl_20575 <= new_AGEMA_signal_3741 & n3665;
  LPM_q_ivl_20578 <= tmp_ivl_20580 & tmp_ivl_20575;
  tmp_ivl_20582 <= tmp_ivl_20586(1);
  tmp_ivl_20584 <= tmp_ivl_20586(0);
  tmp_ivl_20586 <= LPM_d0_ivl_20590(0 + 1 downto 0);
  tmp_ivl_20591 <= new_AGEMA_signal_3589 & n3661;
  LPM_q_ivl_20594 <= tmp_ivl_20596 & tmp_ivl_20591;
  tmp_ivl_20598 <= new_AGEMA_signal_3600 & n3660;
  LPM_q_ivl_20601 <= tmp_ivl_20603 & tmp_ivl_20598;
  new_AGEMA_signal_4017 <= tmp_ivl_20605(1);
  n3662 <= tmp_ivl_20605(0);
  tmp_ivl_20605 <= LPM_d0_ivl_20609(0 + 1 downto 0);
  tmp_ivl_20610 <= new_AGEMA_signal_4017 & n3662;
  LPM_q_ivl_20613 <= tmp_ivl_20615 & tmp_ivl_20610;
  tmp_ivl_20617 <= new_AGEMA_signal_3741 & n3665;
  LPM_q_ivl_20620 <= tmp_ivl_20622 & tmp_ivl_20617;
  tmp_ivl_20624 <= tmp_ivl_20628(1);
  tmp_ivl_20626 <= tmp_ivl_20628(0);
  tmp_ivl_20628 <= LPM_d0_ivl_20632(0 + 1 downto 0);
  tmp_ivl_20633 <= new_AGEMA_signal_3586 & n3664;
  LPM_q_ivl_20636 <= tmp_ivl_20638 & tmp_ivl_20633;
  tmp_ivl_20640 <= new_AGEMA_signal_3588 & n3663;
  LPM_q_ivl_20643 <= tmp_ivl_20645 & tmp_ivl_20640;
  new_AGEMA_signal_4018 <= tmp_ivl_20647(1);
  n3666 <= tmp_ivl_20647(0);
  tmp_ivl_20647 <= LPM_d0_ivl_20651(0 + 1 downto 0);
  tmp_ivl_20652 <= new_AGEMA_signal_4018 & n3666;
  LPM_q_ivl_20655 <= tmp_ivl_20657 & tmp_ivl_20652;
  tmp_ivl_20659 <= new_AGEMA_signal_3741 & n3665;
  LPM_q_ivl_20662 <= tmp_ivl_20664 & tmp_ivl_20659;
  tmp_ivl_20666 <= tmp_ivl_20670(1);
  tmp_ivl_20668 <= tmp_ivl_20670(0);
  tmp_ivl_20670 <= LPM_d0_ivl_20674(0 + 1 downto 0);
  tmp_ivl_20675 <= new_AGEMA_signal_3680 & n3667;
  LPM_q_ivl_20678 <= tmp_ivl_20680 & tmp_ivl_20675;
  tmp_ivl_20682 <= new_AGEMA_signal_3688 & n3863;
  LPM_q_ivl_20685 <= tmp_ivl_20687 & tmp_ivl_20682;
  new_AGEMA_signal_4019 <= tmp_ivl_20689(1);
  n3669 <= tmp_ivl_20689(0);
  tmp_ivl_20689 <= LPM_d0_ivl_20693(0 + 1 downto 0);
  tmp_ivl_20695 <= z0(1);
  tmp_ivl_20696 <= new_AGEMA_signal_3890 & tmp_ivl_20695;
  LPM_q_ivl_20699 <= tmp_ivl_20701 & tmp_ivl_20696;
  tmp_ivl_20704 <= state_in_s1(57);
  tmp_ivl_20706 <= state_in_s0(57);
  tmp_ivl_20707 <= tmp_ivl_20704 & tmp_ivl_20706;
  LPM_q_ivl_20710 <= tmp_ivl_20712 & tmp_ivl_20707;
  new_AGEMA_signal_4020 <= tmp_ivl_20714(1);
  n3673 <= tmp_ivl_20714(0);
  tmp_ivl_20714 <= LPM_d0_ivl_20718(0 + 1 downto 0);
  tmp_ivl_20719 <= new_AGEMA_signal_4020 & n3673;
  LPM_q_ivl_20722 <= tmp_ivl_20724 & tmp_ivl_20719;
  tmp_ivl_20726 <= new_AGEMA_signal_3300 & n3668;
  LPM_q_ivl_20729 <= tmp_ivl_20731 & tmp_ivl_20726;
  new_AGEMA_signal_4319 <= tmp_ivl_20733(1);
  n3842 <= tmp_ivl_20733(0);
  tmp_ivl_20733 <= LPM_d0_ivl_20737(0 + 1 downto 0);
  tmp_ivl_20738 <= new_AGEMA_signal_4019 & n3669;
  LPM_q_ivl_20741 <= tmp_ivl_20743 & tmp_ivl_20738;
  tmp_ivl_20745 <= new_AGEMA_signal_4319 & n3842;
  LPM_q_ivl_20748 <= tmp_ivl_20750 & tmp_ivl_20745;
  tmp_ivl_20752 <= tmp_ivl_20756(1);
  tmp_ivl_20754 <= tmp_ivl_20756(0);
  tmp_ivl_20756 <= LPM_d0_ivl_20760(0 + 1 downto 0);
  tmp_ivl_20761 <= new_AGEMA_signal_3679 & n3671;
  LPM_q_ivl_20764 <= tmp_ivl_20766 & tmp_ivl_20761;
  tmp_ivl_20768 <= new_AGEMA_signal_3706 & n3670;
  LPM_q_ivl_20771 <= tmp_ivl_20773 & tmp_ivl_20768;
  new_AGEMA_signal_4021 <= tmp_ivl_20775(1);
  n3672 <= tmp_ivl_20775(0);
  tmp_ivl_20775 <= LPM_d0_ivl_20779(0 + 1 downto 0);
  tmp_ivl_20780 <= new_AGEMA_signal_4021 & n3672;
  LPM_q_ivl_20783 <= tmp_ivl_20785 & tmp_ivl_20780;
  tmp_ivl_20787 <= new_AGEMA_signal_4319 & n3842;
  LPM_q_ivl_20790 <= tmp_ivl_20792 & tmp_ivl_20787;
  tmp_ivl_20794 <= tmp_ivl_20798(1);
  tmp_ivl_20796 <= tmp_ivl_20798(0);
  tmp_ivl_20798 <= LPM_d0_ivl_20802(0 + 1 downto 0);
  tmp_ivl_20803 <= new_AGEMA_signal_3942 & n3898;
  LPM_q_ivl_20806 <= tmp_ivl_20808 & tmp_ivl_20803;
  tmp_ivl_20810 <= new_AGEMA_signal_3994 & n3790;
  LPM_q_ivl_20813 <= tmp_ivl_20815 & tmp_ivl_20810;
  new_AGEMA_signal_4320 <= tmp_ivl_20817(1);
  n3676 <= tmp_ivl_20817(0);
  tmp_ivl_20817 <= LPM_d0_ivl_20821(0 + 1 downto 0);
  tmp_ivl_20823 <= z1(1);
  tmp_ivl_20824 <= new_AGEMA_signal_3887 & tmp_ivl_20823;
  LPM_q_ivl_20827 <= tmp_ivl_20829 & tmp_ivl_20824;
  tmp_ivl_20832 <= state_in_s1(313);
  tmp_ivl_20834 <= state_in_s0(313);
  tmp_ivl_20835 <= tmp_ivl_20832 & tmp_ivl_20834;
  LPM_q_ivl_20838 <= tmp_ivl_20840 & tmp_ivl_20835;
  new_AGEMA_signal_4022 <= tmp_ivl_20842(1);
  n3675 <= tmp_ivl_20842(0);
  tmp_ivl_20842 <= LPM_d0_ivl_20846(0 + 1 downto 0);
  tmp_ivl_20848 <= state_in_s1(121);
  tmp_ivl_20850 <= state_in_s0(121);
  tmp_ivl_20851 <= tmp_ivl_20848 & tmp_ivl_20850;
  LPM_q_ivl_20854 <= tmp_ivl_20856 & tmp_ivl_20851;
  tmp_ivl_20858 <= new_AGEMA_signal_4020 & n3673;
  LPM_q_ivl_20861 <= tmp_ivl_20863 & tmp_ivl_20858;
  new_AGEMA_signal_4321 <= tmp_ivl_20865(1);
  n3674 <= tmp_ivl_20865(0);
  tmp_ivl_20865 <= LPM_d0_ivl_20869(0 + 1 downto 0);
  tmp_ivl_20870 <= new_AGEMA_signal_4022 & n3675;
  LPM_q_ivl_20873 <= tmp_ivl_20875 & tmp_ivl_20870;
  tmp_ivl_20877 <= new_AGEMA_signal_4321 & n3674;
  LPM_q_ivl_20880 <= tmp_ivl_20882 & tmp_ivl_20877;
  new_AGEMA_signal_4496 <= tmp_ivl_20884(1);
  n3903 <= tmp_ivl_20884(0);
  tmp_ivl_20884 <= LPM_d0_ivl_20888(0 + 1 downto 0);
  tmp_ivl_20889 <= new_AGEMA_signal_4320 & n3676;
  LPM_q_ivl_20892 <= tmp_ivl_20894 & tmp_ivl_20889;
  tmp_ivl_20896 <= new_AGEMA_signal_4496 & n3903;
  LPM_q_ivl_20899 <= tmp_ivl_20901 & tmp_ivl_20896;
  tmp_ivl_20903 <= tmp_ivl_20907(1);
  tmp_ivl_20905 <= tmp_ivl_20907(0);
  tmp_ivl_20907 <= LPM_d0_ivl_20911(0 + 1 downto 0);
  tmp_ivl_20912 <= new_AGEMA_signal_3988 & n3678;
  LPM_q_ivl_20915 <= tmp_ivl_20917 & tmp_ivl_20912;
  tmp_ivl_20919 <= new_AGEMA_signal_3993 & n3677;
  LPM_q_ivl_20922 <= tmp_ivl_20924 & tmp_ivl_20919;
  new_AGEMA_signal_4322 <= tmp_ivl_20926(1);
  n3679 <= tmp_ivl_20926(0);
  tmp_ivl_20926 <= LPM_d0_ivl_20930(0 + 1 downto 0);
  tmp_ivl_20931 <= new_AGEMA_signal_4322 & n3679;
  LPM_q_ivl_20934 <= tmp_ivl_20936 & tmp_ivl_20931;
  tmp_ivl_20938 <= new_AGEMA_signal_4496 & n3903;
  LPM_q_ivl_20941 <= tmp_ivl_20943 & tmp_ivl_20938;
  tmp_ivl_20945 <= tmp_ivl_20949(1);
  tmp_ivl_20947 <= tmp_ivl_20949(0);
  tmp_ivl_20949 <= LPM_d0_ivl_20953(0 + 1 downto 0);
  tmp_ivl_20954 <= new_AGEMA_signal_3425 & n3681;
  LPM_q_ivl_20957 <= tmp_ivl_20959 & tmp_ivl_20954;
  tmp_ivl_20961 <= new_AGEMA_signal_3403 & n3680;
  LPM_q_ivl_20964 <= tmp_ivl_20966 & tmp_ivl_20961;
  new_AGEMA_signal_3742 <= tmp_ivl_20968(1);
  n3914 <= tmp_ivl_20968(0);
  tmp_ivl_20968 <= LPM_d0_ivl_20972(0 + 1 downto 0);
  tmp_ivl_20974 <= state_in_s1(232);
  tmp_ivl_20976 <= state_in_s0(232);
  tmp_ivl_20977 <= tmp_ivl_20974 & tmp_ivl_20976;
  LPM_q_ivl_20980 <= tmp_ivl_20982 & tmp_ivl_20977;
  tmp_ivl_20985 <= z4(16);
  tmp_ivl_20986 <= new_AGEMA_signal_3118 & tmp_ivl_20985;
  LPM_q_ivl_20989 <= tmp_ivl_20991 & tmp_ivl_20986;
  new_AGEMA_signal_3444 <= tmp_ivl_20993(1);
  n3688 <= tmp_ivl_20993(0);
  tmp_ivl_20993 <= LPM_d0_ivl_20997(0 + 1 downto 0);
  tmp_ivl_20998 <= new_AGEMA_signal_3357 & n3682;
  LPM_q_ivl_21001 <= tmp_ivl_21003 & tmp_ivl_20998;
  tmp_ivl_21005 <= new_AGEMA_signal_3444 & n3688;
  LPM_q_ivl_21008 <= tmp_ivl_21010 & tmp_ivl_21005;
  new_AGEMA_signal_3743 <= tmp_ivl_21012(1);
  n3911 <= tmp_ivl_21012(0);
  tmp_ivl_21012 <= LPM_d0_ivl_21016(0 + 1 downto 0);
  tmp_ivl_21017 <= new_AGEMA_signal_3742 & n3914;
  LPM_q_ivl_21020 <= tmp_ivl_21022 & tmp_ivl_21017;
  tmp_ivl_21024 <= new_AGEMA_signal_3743 & n3911;
  LPM_q_ivl_21027 <= tmp_ivl_21029 & tmp_ivl_21024;
  new_AGEMA_signal_4023 <= tmp_ivl_21031(1);
  n3685 <= tmp_ivl_21031(0);
  tmp_ivl_21031 <= LPM_d0_ivl_21035(0 + 1 downto 0);
  tmp_ivl_21036 <= new_AGEMA_signal_3372 & n3684;
  LPM_q_ivl_21039 <= tmp_ivl_21041 & tmp_ivl_21036;
  tmp_ivl_21043 <= new_AGEMA_signal_3365 & n3683;
  LPM_q_ivl_21046 <= tmp_ivl_21048 & tmp_ivl_21043;
  new_AGEMA_signal_3744 <= tmp_ivl_21050(1);
  n3759 <= tmp_ivl_21050(0);
  tmp_ivl_21050 <= LPM_d0_ivl_21054(0 + 1 downto 0);
  tmp_ivl_21055 <= new_AGEMA_signal_4023 & n3685;
  LPM_q_ivl_21058 <= tmp_ivl_21060 & tmp_ivl_21055;
  tmp_ivl_21062 <= new_AGEMA_signal_3744 & n3759;
  LPM_q_ivl_21065 <= tmp_ivl_21067 & tmp_ivl_21062;
  tmp_ivl_21069 <= tmp_ivl_21073(1);
  tmp_ivl_21071 <= tmp_ivl_21073(0);
  tmp_ivl_21073 <= LPM_d0_ivl_21077(0 + 1 downto 0);
  tmp_ivl_21078 <= new_AGEMA_signal_3603 & n3687;
  LPM_q_ivl_21081 <= tmp_ivl_21083 & tmp_ivl_21078;
  tmp_ivl_21085 <= new_AGEMA_signal_3610 & n3686;
  LPM_q_ivl_21088 <= tmp_ivl_21090 & tmp_ivl_21085;
  new_AGEMA_signal_4024 <= tmp_ivl_21092(1);
  n3689 <= tmp_ivl_21092(0);
  tmp_ivl_21092 <= LPM_d0_ivl_21096(0 + 1 downto 0);
  tmp_ivl_21098 <= state_in_s1(296);
  tmp_ivl_21100 <= state_in_s0(296);
  tmp_ivl_21101 <= tmp_ivl_21098 & tmp_ivl_21100;
  LPM_q_ivl_21104 <= tmp_ivl_21106 & tmp_ivl_21101;
  tmp_ivl_21108 <= new_AGEMA_signal_3444 & n3688;
  LPM_q_ivl_21111 <= tmp_ivl_21113 & tmp_ivl_21108;
  new_AGEMA_signal_3745 <= tmp_ivl_21115(1);
  n3732 <= tmp_ivl_21115(0);
  tmp_ivl_21115 <= LPM_d0_ivl_21119(0 + 1 downto 0);
  tmp_ivl_21120 <= new_AGEMA_signal_4024 & n3689;
  LPM_q_ivl_21123 <= tmp_ivl_21125 & tmp_ivl_21120;
  tmp_ivl_21127 <= new_AGEMA_signal_3745 & n3732;
  LPM_q_ivl_21130 <= tmp_ivl_21132 & tmp_ivl_21127;
  tmp_ivl_21134 <= tmp_ivl_21138(1);
  tmp_ivl_21136 <= tmp_ivl_21138(0);
  tmp_ivl_21138 <= LPM_d0_ivl_21142(0 + 1 downto 0);
  tmp_ivl_21143 <= new_AGEMA_signal_3630 & n3726;
  LPM_q_ivl_21146 <= tmp_ivl_21148 & tmp_ivl_21143;
  tmp_ivl_21150 <= new_AGEMA_signal_3727 & n3690;
  LPM_q_ivl_21153 <= tmp_ivl_21155 & tmp_ivl_21150;
  new_AGEMA_signal_4025 <= tmp_ivl_21157(1);
  n3691 <= tmp_ivl_21157(0);
  tmp_ivl_21157 <= LPM_d0_ivl_21161(0 + 1 downto 0);
  tmp_ivl_21162 <= new_AGEMA_signal_4025 & n3691;
  LPM_q_ivl_21165 <= tmp_ivl_21167 & tmp_ivl_21162;
  tmp_ivl_21169 <= new_AGEMA_signal_3745 & n3732;
  LPM_q_ivl_21172 <= tmp_ivl_21174 & tmp_ivl_21169;
  tmp_ivl_21176 <= tmp_ivl_21180(1);
  tmp_ivl_21178 <= tmp_ivl_21180(0);
  tmp_ivl_21180 <= LPM_d0_ivl_21184(0 + 1 downto 0);
  tmp_ivl_21185 <= new_AGEMA_signal_3673 & n3774;
  LPM_q_ivl_21188 <= tmp_ivl_21190 & tmp_ivl_21185;
  tmp_ivl_21192 <= new_AGEMA_signal_3721 & n3855;
  LPM_q_ivl_21195 <= tmp_ivl_21197 & tmp_ivl_21192;
  new_AGEMA_signal_4026 <= tmp_ivl_21199(1);
  n3693 <= tmp_ivl_21199(0);
  tmp_ivl_21199 <= LPM_d0_ivl_21203(0 + 1 downto 0);
  tmp_ivl_21205 <= z0(44);
  tmp_ivl_21206 <= new_AGEMA_signal_3215 & tmp_ivl_21205;
  LPM_q_ivl_21209 <= tmp_ivl_21211 & tmp_ivl_21206;
  tmp_ivl_21214 <= state_in_s1(20);
  tmp_ivl_21216 <= state_in_s0(20);
  tmp_ivl_21217 <= tmp_ivl_21214 & tmp_ivl_21216;
  LPM_q_ivl_21220 <= tmp_ivl_21222 & tmp_ivl_21217;
  new_AGEMA_signal_3445 <= tmp_ivl_21224(1);
  n3698 <= tmp_ivl_21224(0);
  tmp_ivl_21224 <= LPM_d0_ivl_21228(0 + 1 downto 0);
  tmp_ivl_21229 <= new_AGEMA_signal_3445 & n3698;
  LPM_q_ivl_21232 <= tmp_ivl_21234 & tmp_ivl_21229;
  tmp_ivl_21236 <= new_AGEMA_signal_3305 & n3692;
  LPM_q_ivl_21239 <= tmp_ivl_21241 & tmp_ivl_21236;
  new_AGEMA_signal_3746 <= tmp_ivl_21243(1);
  n3695 <= tmp_ivl_21243(0);
  tmp_ivl_21243 <= LPM_d0_ivl_21247(0 + 1 downto 0);
  tmp_ivl_21248 <= new_AGEMA_signal_4026 & n3693;
  LPM_q_ivl_21251 <= tmp_ivl_21253 & tmp_ivl_21248;
  tmp_ivl_21255 <= new_AGEMA_signal_3746 & n3695;
  LPM_q_ivl_21258 <= tmp_ivl_21260 & tmp_ivl_21255;
  tmp_ivl_21262 <= tmp_ivl_21266(1);
  tmp_ivl_21264 <= tmp_ivl_21266(0);
  tmp_ivl_21266 <= LPM_d0_ivl_21270(0 + 1 downto 0);
  tmp_ivl_21271 <= new_AGEMA_signal_3715 & n3773;
  LPM_q_ivl_21274 <= tmp_ivl_21276 & tmp_ivl_21271;
  tmp_ivl_21278 <= new_AGEMA_signal_3744 & n3759;
  LPM_q_ivl_21281 <= tmp_ivl_21283 & tmp_ivl_21278;
  new_AGEMA_signal_4027 <= tmp_ivl_21285(1);
  n3694 <= tmp_ivl_21285(0);
  tmp_ivl_21285 <= LPM_d0_ivl_21289(0 + 1 downto 0);
  tmp_ivl_21290 <= new_AGEMA_signal_4027 & n3694;
  LPM_q_ivl_21293 <= tmp_ivl_21295 & tmp_ivl_21290;
  tmp_ivl_21297 <= new_AGEMA_signal_3746 & n3695;
  LPM_q_ivl_21300 <= tmp_ivl_21302 & tmp_ivl_21297;
  tmp_ivl_21304 <= tmp_ivl_21308(1);
  tmp_ivl_21306 <= tmp_ivl_21308(0);
  tmp_ivl_21308 <= LPM_d0_ivl_21312(0 + 1 downto 0);
  tmp_ivl_21313 <= new_AGEMA_signal_3719 & n3876;
  LPM_q_ivl_21316 <= tmp_ivl_21318 & tmp_ivl_21313;
  tmp_ivl_21320 <= new_AGEMA_signal_3743 & n3911;
  LPM_q_ivl_21323 <= tmp_ivl_21325 & tmp_ivl_21320;
  new_AGEMA_signal_4028 <= tmp_ivl_21327(1);
  n3696 <= tmp_ivl_21327(0);
  tmp_ivl_21327 <= LPM_d0_ivl_21331(0 + 1 downto 0);
  tmp_ivl_21332 <= new_AGEMA_signal_4028 & n3696;
  LPM_q_ivl_21335 <= tmp_ivl_21337 & tmp_ivl_21332;
  tmp_ivl_21339 <= new_AGEMA_signal_3746 & n3695;
  LPM_q_ivl_21342 <= tmp_ivl_21344 & tmp_ivl_21339;
  tmp_ivl_21346 <= tmp_ivl_21350(1);
  tmp_ivl_21348 <= tmp_ivl_21350(0);
  tmp_ivl_21350 <= LPM_d0_ivl_21354(0 + 1 downto 0);
  tmp_ivl_21355 <= new_AGEMA_signal_3921 & n3697;
  LPM_q_ivl_21358 <= tmp_ivl_21360 & tmp_ivl_21355;
  tmp_ivl_21362 <= new_AGEMA_signal_4001 & n3719;
  LPM_q_ivl_21365 <= tmp_ivl_21367 & tmp_ivl_21362;
  new_AGEMA_signal_4329 <= tmp_ivl_21369(1);
  n3701 <= tmp_ivl_21369(0);
  tmp_ivl_21369 <= LPM_d0_ivl_21373(0 + 1 downto 0);
  tmp_ivl_21375 <= z1(44);
  tmp_ivl_21376 <= new_AGEMA_signal_3025 & tmp_ivl_21375;
  LPM_q_ivl_21379 <= tmp_ivl_21381 & tmp_ivl_21376;
  tmp_ivl_21383 <= new_AGEMA_signal_3445 & n3698;
  LPM_q_ivl_21386 <= tmp_ivl_21388 & tmp_ivl_21383;
  new_AGEMA_signal_3747 <= tmp_ivl_21390(1);
  n3700 <= tmp_ivl_21390(0);
  tmp_ivl_21390 <= LPM_d0_ivl_21394(0 + 1 downto 0);
  tmp_ivl_21395 <= new_AGEMA_signal_3747 & n3700;
  LPM_q_ivl_21398 <= tmp_ivl_21400 & tmp_ivl_21395;
  tmp_ivl_21402 <= new_AGEMA_signal_2687 & n3699;
  LPM_q_ivl_21405 <= tmp_ivl_21407 & tmp_ivl_21402;
  new_AGEMA_signal_4029 <= tmp_ivl_21409(1);
  n3754 <= tmp_ivl_21409(0);
  tmp_ivl_21409 <= LPM_d0_ivl_21413(0 + 1 downto 0);
  tmp_ivl_21414 <= new_AGEMA_signal_4329 & n3701;
  LPM_q_ivl_21417 <= tmp_ivl_21419 & tmp_ivl_21414;
  tmp_ivl_21421 <= new_AGEMA_signal_4029 & n3754;
  LPM_q_ivl_21424 <= tmp_ivl_21426 & tmp_ivl_21421;
  tmp_ivl_21428 <= tmp_ivl_21432(1);
  tmp_ivl_21430 <= tmp_ivl_21432(0);
  tmp_ivl_21432 <= LPM_d0_ivl_21436(0 + 1 downto 0);
  tmp_ivl_21437 <= new_AGEMA_signal_3935 & n3750;
  LPM_q_ivl_21440 <= tmp_ivl_21442 & tmp_ivl_21437;
  tmp_ivl_21444 <= new_AGEMA_signal_3986 & n3702;
  LPM_q_ivl_21447 <= tmp_ivl_21449 & tmp_ivl_21444;
  new_AGEMA_signal_4330 <= tmp_ivl_21451(1);
  n3703 <= tmp_ivl_21451(0);
  tmp_ivl_21451 <= LPM_d0_ivl_21455(0 + 1 downto 0);
  tmp_ivl_21456 <= new_AGEMA_signal_4330 & n3703;
  LPM_q_ivl_21459 <= tmp_ivl_21461 & tmp_ivl_21456;
  tmp_ivl_21463 <= new_AGEMA_signal_4029 & n3754;
  LPM_q_ivl_21466 <= tmp_ivl_21468 & tmp_ivl_21463;
  tmp_ivl_21470 <= tmp_ivl_21474(1);
  tmp_ivl_21472 <= tmp_ivl_21474(0);
  tmp_ivl_21474 <= LPM_d0_ivl_21478(0 + 1 downto 0);
  tmp_ivl_21479 <= new_AGEMA_signal_3644 & n3705;
  LPM_q_ivl_21482 <= tmp_ivl_21484 & tmp_ivl_21479;
  tmp_ivl_21486 <= new_AGEMA_signal_3678 & n3704;
  LPM_q_ivl_21489 <= tmp_ivl_21491 & tmp_ivl_21486;
  new_AGEMA_signal_4030 <= tmp_ivl_21493(1);
  n3707 <= tmp_ivl_21493(0);
  tmp_ivl_21493 <= LPM_d0_ivl_21497(0 + 1 downto 0);
  tmp_ivl_21499 <= z0(2);
  tmp_ivl_21500 <= new_AGEMA_signal_4203 & tmp_ivl_21499;
  LPM_q_ivl_21503 <= tmp_ivl_21505 & tmp_ivl_21500;
  tmp_ivl_21508 <= state_in_s1(58);
  tmp_ivl_21510 <= state_in_s0(58);
  tmp_ivl_21511 <= tmp_ivl_21508 & tmp_ivl_21510;
  LPM_q_ivl_21514 <= tmp_ivl_21516 & tmp_ivl_21511;
  new_AGEMA_signal_4331 <= tmp_ivl_21518(1);
  n3715 <= tmp_ivl_21518(0);
  tmp_ivl_21518 <= LPM_d0_ivl_21522(0 + 1 downto 0);
  tmp_ivl_21523 <= new_AGEMA_signal_4331 & n3715;
  LPM_q_ivl_21526 <= tmp_ivl_21528 & tmp_ivl_21523;
  tmp_ivl_21530 <= new_AGEMA_signal_3303 & n3706;
  LPM_q_ivl_21533 <= tmp_ivl_21535 & tmp_ivl_21530;
  new_AGEMA_signal_4499 <= tmp_ivl_21537(1);
  n3713 <= tmp_ivl_21537(0);
  tmp_ivl_21537 <= LPM_d0_ivl_21541(0 + 1 downto 0);
  tmp_ivl_21542 <= new_AGEMA_signal_4030 & n3707;
  LPM_q_ivl_21545 <= tmp_ivl_21547 & tmp_ivl_21542;
  tmp_ivl_21549 <= new_AGEMA_signal_4499 & n3713;
  LPM_q_ivl_21552 <= tmp_ivl_21554 & tmp_ivl_21549;
  tmp_ivl_21556 <= tmp_ivl_21560(1);
  tmp_ivl_21558 <= tmp_ivl_21560(0);
  tmp_ivl_21560 <= LPM_d0_ivl_21564(0 + 1 downto 0);
  tmp_ivl_21565 <= new_AGEMA_signal_3643 & n3709;
  LPM_q_ivl_21568 <= tmp_ivl_21570 & tmp_ivl_21565;
  tmp_ivl_21572 <= new_AGEMA_signal_3697 & n3708;
  LPM_q_ivl_21575 <= tmp_ivl_21577 & tmp_ivl_21572;
  new_AGEMA_signal_4031 <= tmp_ivl_21579(1);
  n3710 <= tmp_ivl_21579(0);
  tmp_ivl_21579 <= LPM_d0_ivl_21583(0 + 1 downto 0);
  tmp_ivl_21584 <= new_AGEMA_signal_4031 & n3710;
  LPM_q_ivl_21587 <= tmp_ivl_21589 & tmp_ivl_21584;
  tmp_ivl_21591 <= new_AGEMA_signal_4499 & n3713;
  LPM_q_ivl_21594 <= tmp_ivl_21596 & tmp_ivl_21591;
  tmp_ivl_21598 <= tmp_ivl_21602(1);
  tmp_ivl_21600 <= tmp_ivl_21602(0);
  tmp_ivl_21602 <= LPM_d0_ivl_21606(0 + 1 downto 0);
  tmp_ivl_21607 <= new_AGEMA_signal_3696 & n3712;
  LPM_q_ivl_21610 <= tmp_ivl_21612 & tmp_ivl_21607;
  tmp_ivl_21614 <= new_AGEMA_signal_3734 & n3711;
  LPM_q_ivl_21617 <= tmp_ivl_21619 & tmp_ivl_21614;
  new_AGEMA_signal_4032 <= tmp_ivl_21621(1);
  n3714 <= tmp_ivl_21621(0);
  tmp_ivl_21621 <= LPM_d0_ivl_21625(0 + 1 downto 0);
  tmp_ivl_21626 <= new_AGEMA_signal_4032 & n3714;
  LPM_q_ivl_21629 <= tmp_ivl_21631 & tmp_ivl_21626;
  tmp_ivl_21633 <= new_AGEMA_signal_4499 & n3713;
  LPM_q_ivl_21636 <= tmp_ivl_21638 & tmp_ivl_21633;
  tmp_ivl_21640 <= tmp_ivl_21644(1);
  tmp_ivl_21642 <= tmp_ivl_21644(0);
  tmp_ivl_21644 <= LPM_d0_ivl_21648(0 + 1 downto 0);
  tmp_ivl_21649 <= new_AGEMA_signal_3956 & n3744;
  LPM_q_ivl_21652 <= tmp_ivl_21654 & tmp_ivl_21649;
  tmp_ivl_21656 <= new_AGEMA_signal_3997 & n3848;
  LPM_q_ivl_21659 <= tmp_ivl_21661 & tmp_ivl_21656;
  new_AGEMA_signal_4332 <= tmp_ivl_21663(1);
  n3718 <= tmp_ivl_21663(0);
  tmp_ivl_21663 <= LPM_d0_ivl_21667(0 + 1 downto 0);
  tmp_ivl_21669 <= z1(2);
  tmp_ivl_21670 <= new_AGEMA_signal_4200 & tmp_ivl_21669;
  LPM_q_ivl_21673 <= tmp_ivl_21675 & tmp_ivl_21670;
  tmp_ivl_21678 <= state_in_s1(314);
  tmp_ivl_21680 <= state_in_s0(314);
  tmp_ivl_21681 <= tmp_ivl_21678 & tmp_ivl_21680;
  LPM_q_ivl_21684 <= tmp_ivl_21686 & tmp_ivl_21681;
  new_AGEMA_signal_4333 <= tmp_ivl_21688(1);
  n3717 <= tmp_ivl_21688(0);
  tmp_ivl_21688 <= LPM_d0_ivl_21692(0 + 1 downto 0);
  tmp_ivl_21694 <= state_in_s1(122);
  tmp_ivl_21696 <= state_in_s0(122);
  tmp_ivl_21697 <= tmp_ivl_21694 & tmp_ivl_21696;
  LPM_q_ivl_21700 <= tmp_ivl_21702 & tmp_ivl_21697;
  tmp_ivl_21704 <= new_AGEMA_signal_4331 & n3715;
  LPM_q_ivl_21707 <= tmp_ivl_21709 & tmp_ivl_21704;
  new_AGEMA_signal_4500 <= tmp_ivl_21711(1);
  n3716 <= tmp_ivl_21711(0);
  tmp_ivl_21711 <= LPM_d0_ivl_21715(0 + 1 downto 0);
  tmp_ivl_21716 <= new_AGEMA_signal_4333 & n3717;
  LPM_q_ivl_21719 <= tmp_ivl_21721 & tmp_ivl_21716;
  tmp_ivl_21723 <= new_AGEMA_signal_4500 & n3716;
  LPM_q_ivl_21726 <= tmp_ivl_21728 & tmp_ivl_21723;
  new_AGEMA_signal_4586 <= tmp_ivl_21730(1);
  n3753 <= tmp_ivl_21730(0);
  tmp_ivl_21730 <= LPM_d0_ivl_21734(0 + 1 downto 0);
  tmp_ivl_21735 <= new_AGEMA_signal_4332 & n3718;
  LPM_q_ivl_21738 <= tmp_ivl_21740 & tmp_ivl_21735;
  tmp_ivl_21742 <= new_AGEMA_signal_4586 & n3753;
  LPM_q_ivl_21745 <= tmp_ivl_21747 & tmp_ivl_21742;
  tmp_ivl_21749 <= tmp_ivl_21753(1);
  tmp_ivl_21751 <= tmp_ivl_21753(0);
  tmp_ivl_21753 <= LPM_d0_ivl_21757(0 + 1 downto 0);
  tmp_ivl_21758 <= new_AGEMA_signal_3996 & n3720;
  LPM_q_ivl_21761 <= tmp_ivl_21763 & tmp_ivl_21758;
  tmp_ivl_21765 <= new_AGEMA_signal_4001 & n3719;
  LPM_q_ivl_21768 <= tmp_ivl_21770 & tmp_ivl_21765;
  new_AGEMA_signal_4334 <= tmp_ivl_21772(1);
  n3721 <= tmp_ivl_21772(0);
  tmp_ivl_21772 <= LPM_d0_ivl_21776(0 + 1 downto 0);
  tmp_ivl_21777 <= new_AGEMA_signal_4334 & n3721;
  LPM_q_ivl_21780 <= tmp_ivl_21782 & tmp_ivl_21777;
  tmp_ivl_21784 <= new_AGEMA_signal_4586 & n3753;
  LPM_q_ivl_21787 <= tmp_ivl_21789 & tmp_ivl_21784;
  tmp_ivl_21791 <= tmp_ivl_21795(1);
  tmp_ivl_21793 <= tmp_ivl_21795(0);
  tmp_ivl_21795 <= LPM_d0_ivl_21799(0 + 1 downto 0);
  tmp_ivl_21800 <= new_AGEMA_signal_3711 & n3805;
  LPM_q_ivl_21803 <= tmp_ivl_21805 & tmp_ivl_21800;
  tmp_ivl_21807 <= new_AGEMA_signal_3725 & n3890;
  LPM_q_ivl_21810 <= tmp_ivl_21812 & tmp_ivl_21807;
  new_AGEMA_signal_4033 <= tmp_ivl_21814(1);
  n3723 <= tmp_ivl_21814(0);
  tmp_ivl_21814 <= LPM_d0_ivl_21818(0 + 1 downto 0);
  tmp_ivl_21820 <= state_in_s1(202);
  tmp_ivl_21822 <= state_in_s0(202);
  tmp_ivl_21823 <= tmp_ivl_21820 & tmp_ivl_21822;
  LPM_q_ivl_21826 <= tmp_ivl_21828 & tmp_ivl_21823;
  tmp_ivl_21831 <= z4(50);
  tmp_ivl_21832 <= new_AGEMA_signal_3156 & tmp_ivl_21831;
  LPM_q_ivl_21835 <= tmp_ivl_21837 & tmp_ivl_21832;
  new_AGEMA_signal_3446 <= tmp_ivl_21839(1);
  n3727 <= tmp_ivl_21839(0);
  tmp_ivl_21839 <= LPM_d0_ivl_21843(0 + 1 downto 0);
  tmp_ivl_21844 <= new_AGEMA_signal_3374 & n3722;
  LPM_q_ivl_21847 <= tmp_ivl_21849 & tmp_ivl_21844;
  tmp_ivl_21851 <= new_AGEMA_signal_3446 & n3727;
  LPM_q_ivl_21854 <= tmp_ivl_21856 & tmp_ivl_21851;
  new_AGEMA_signal_3748 <= tmp_ivl_21858(1);
  n3736 <= tmp_ivl_21858(0);
  tmp_ivl_21858 <= LPM_d0_ivl_21862(0 + 1 downto 0);
  tmp_ivl_21863 <= new_AGEMA_signal_4033 & n3723;
  LPM_q_ivl_21866 <= tmp_ivl_21868 & tmp_ivl_21863;
  tmp_ivl_21870 <= new_AGEMA_signal_3748 & n3736;
  LPM_q_ivl_21873 <= tmp_ivl_21875 & tmp_ivl_21870;
  tmp_ivl_21877 <= tmp_ivl_21881(1);
  tmp_ivl_21879 <= tmp_ivl_21881(0);
  tmp_ivl_21881 <= LPM_d0_ivl_21885(0 + 1 downto 0);
  tmp_ivl_21886 <= new_AGEMA_signal_3667 & n3806;
  LPM_q_ivl_21889 <= tmp_ivl_21891 & tmp_ivl_21886;
  tmp_ivl_21893 <= new_AGEMA_signal_3729 & n3740;
  LPM_q_ivl_21896 <= tmp_ivl_21898 & tmp_ivl_21893;
  new_AGEMA_signal_4034 <= tmp_ivl_21900(1);
  n3724 <= tmp_ivl_21900(0);
  tmp_ivl_21900 <= LPM_d0_ivl_21904(0 + 1 downto 0);
  tmp_ivl_21905 <= new_AGEMA_signal_4034 & n3724;
  LPM_q_ivl_21908 <= tmp_ivl_21910 & tmp_ivl_21905;
  tmp_ivl_21912 <= new_AGEMA_signal_3748 & n3736;
  LPM_q_ivl_21915 <= tmp_ivl_21917 & tmp_ivl_21912;
  tmp_ivl_21919 <= tmp_ivl_21923(1);
  tmp_ivl_21921 <= tmp_ivl_21923(0);
  tmp_ivl_21923 <= LPM_d0_ivl_21927(0 + 1 downto 0);
  tmp_ivl_21928 <= new_AGEMA_signal_3630 & n3726;
  LPM_q_ivl_21931 <= tmp_ivl_21933 & tmp_ivl_21928;
  tmp_ivl_21935 <= new_AGEMA_signal_3674 & n3725;
  LPM_q_ivl_21938 <= tmp_ivl_21940 & tmp_ivl_21935;
  new_AGEMA_signal_4035 <= tmp_ivl_21942(1);
  n3728 <= tmp_ivl_21942(0);
  tmp_ivl_21942 <= LPM_d0_ivl_21946(0 + 1 downto 0);
  tmp_ivl_21948 <= state_in_s1(266);
  tmp_ivl_21950 <= state_in_s0(266);
  tmp_ivl_21951 <= tmp_ivl_21948 & tmp_ivl_21950;
  LPM_q_ivl_21954 <= tmp_ivl_21956 & tmp_ivl_21951;
  tmp_ivl_21958 <= new_AGEMA_signal_3446 & n3727;
  LPM_q_ivl_21961 <= tmp_ivl_21963 & tmp_ivl_21958;
  new_AGEMA_signal_3749 <= tmp_ivl_21965(1);
  n3734 <= tmp_ivl_21965(0);
  tmp_ivl_21965 <= LPM_d0_ivl_21969(0 + 1 downto 0);
  tmp_ivl_21970 <= new_AGEMA_signal_4035 & n3728;
  LPM_q_ivl_21973 <= tmp_ivl_21975 & tmp_ivl_21970;
  tmp_ivl_21977 <= new_AGEMA_signal_3749 & n3734;
  LPM_q_ivl_21980 <= tmp_ivl_21982 & tmp_ivl_21977;
  tmp_ivl_21984 <= tmp_ivl_21988(1);
  tmp_ivl_21986 <= tmp_ivl_21988(0);
  tmp_ivl_21988 <= LPM_d0_ivl_21992(0 + 1 downto 0);
  tmp_ivl_21993 <= new_AGEMA_signal_3592 & n3730;
  LPM_q_ivl_21996 <= tmp_ivl_21998 & tmp_ivl_21993;
  tmp_ivl_22000 <= new_AGEMA_signal_3605 & n3729;
  LPM_q_ivl_22003 <= tmp_ivl_22005 & tmp_ivl_22000;
  new_AGEMA_signal_4036 <= tmp_ivl_22007(1);
  n3731 <= tmp_ivl_22007(0);
  tmp_ivl_22007 <= LPM_d0_ivl_22011(0 + 1 downto 0);
  tmp_ivl_22012 <= new_AGEMA_signal_4036 & n3731;
  LPM_q_ivl_22015 <= tmp_ivl_22017 & tmp_ivl_22012;
  tmp_ivl_22019 <= new_AGEMA_signal_3749 & n3734;
  LPM_q_ivl_22022 <= tmp_ivl_22024 & tmp_ivl_22019;
  tmp_ivl_22026 <= tmp_ivl_22030(1);
  tmp_ivl_22028 <= tmp_ivl_22030(0);
  tmp_ivl_22030 <= LPM_d0_ivl_22034(0 + 1 downto 0);
  tmp_ivl_22035 <= new_AGEMA_signal_3591 & n3733;
  LPM_q_ivl_22038 <= tmp_ivl_22040 & tmp_ivl_22035;
  tmp_ivl_22042 <= new_AGEMA_signal_3745 & n3732;
  LPM_q_ivl_22045 <= tmp_ivl_22047 & tmp_ivl_22042;
  new_AGEMA_signal_4037 <= tmp_ivl_22049(1);
  n3735 <= tmp_ivl_22049(0);
  tmp_ivl_22049 <= LPM_d0_ivl_22053(0 + 1 downto 0);
  tmp_ivl_22054 <= new_AGEMA_signal_4037 & n3735;
  LPM_q_ivl_22057 <= tmp_ivl_22059 & tmp_ivl_22054;
  tmp_ivl_22061 <= new_AGEMA_signal_3749 & n3734;
  LPM_q_ivl_22064 <= tmp_ivl_22066 & tmp_ivl_22061;
  tmp_ivl_22068 <= tmp_ivl_22072(1);
  tmp_ivl_22070 <= tmp_ivl_22072(0);
  tmp_ivl_22072 <= LPM_d0_ivl_22076(0 + 1 downto 0);
  tmp_ivl_22077 <= new_AGEMA_signal_3726 & n3737;
  LPM_q_ivl_22080 <= tmp_ivl_22082 & tmp_ivl_22077;
  tmp_ivl_22084 <= new_AGEMA_signal_3748 & n3736;
  LPM_q_ivl_22087 <= tmp_ivl_22089 & tmp_ivl_22084;
  new_AGEMA_signal_4038 <= tmp_ivl_22091(1);
  n3739 <= tmp_ivl_22091(0);
  tmp_ivl_22091 <= LPM_d0_ivl_22095(0 + 1 downto 0);
  tmp_ivl_22097 <= z0(5);
  tmp_ivl_22098 <= new_AGEMA_signal_3889 & tmp_ivl_22097;
  LPM_q_ivl_22101 <= tmp_ivl_22103 & tmp_ivl_22098;
  tmp_ivl_22106 <= state_in_s1(61);
  tmp_ivl_22108 <= state_in_s0(61);
  tmp_ivl_22109 <= tmp_ivl_22106 & tmp_ivl_22108;
  LPM_q_ivl_22112 <= tmp_ivl_22114 & tmp_ivl_22109;
  new_AGEMA_signal_4039 <= tmp_ivl_22116(1);
  n3746 <= tmp_ivl_22116(0);
  tmp_ivl_22116 <= LPM_d0_ivl_22120(0 + 1 downto 0);
  tmp_ivl_22121 <= new_AGEMA_signal_4039 & n3746;
  LPM_q_ivl_22124 <= tmp_ivl_22126 & tmp_ivl_22121;
  tmp_ivl_22128 <= new_AGEMA_signal_3314 & n3738;
  LPM_q_ivl_22131 <= tmp_ivl_22133 & tmp_ivl_22128;
  new_AGEMA_signal_4340 <= tmp_ivl_22135(1);
  n3742 <= tmp_ivl_22135(0);
  tmp_ivl_22135 <= LPM_d0_ivl_22139(0 + 1 downto 0);
  tmp_ivl_22140 <= new_AGEMA_signal_4038 & n3739;
  LPM_q_ivl_22143 <= tmp_ivl_22145 & tmp_ivl_22140;
  tmp_ivl_22147 <= new_AGEMA_signal_4340 & n3742;
  LPM_q_ivl_22150 <= tmp_ivl_22152 & tmp_ivl_22147;
  tmp_ivl_22154 <= tmp_ivl_22158(1);
  tmp_ivl_22156 <= tmp_ivl_22158(0);
  tmp_ivl_22158 <= LPM_d0_ivl_22162(0 + 1 downto 0);
  tmp_ivl_22163 <= new_AGEMA_signal_3692 & n3826;
  LPM_q_ivl_22166 <= tmp_ivl_22168 & tmp_ivl_22163;
  tmp_ivl_22170 <= new_AGEMA_signal_3729 & n3740;
  LPM_q_ivl_22173 <= tmp_ivl_22175 & tmp_ivl_22170;
  new_AGEMA_signal_4040 <= tmp_ivl_22177(1);
  n3741 <= tmp_ivl_22177(0);
  tmp_ivl_22177 <= LPM_d0_ivl_22181(0 + 1 downto 0);
  tmp_ivl_22182 <= new_AGEMA_signal_4040 & n3741;
  LPM_q_ivl_22185 <= tmp_ivl_22187 & tmp_ivl_22182;
  tmp_ivl_22189 <= new_AGEMA_signal_4340 & n3742;
  LPM_q_ivl_22192 <= tmp_ivl_22194 & tmp_ivl_22189;
  tmp_ivl_22196 <= tmp_ivl_22200(1);
  tmp_ivl_22198 <= tmp_ivl_22200(0);
  tmp_ivl_22200 <= LPM_d0_ivl_22204(0 + 1 downto 0);
  tmp_ivl_22205 <= new_AGEMA_signal_3691 & n3918;
  LPM_q_ivl_22208 <= tmp_ivl_22210 & tmp_ivl_22205;
  tmp_ivl_22212 <= new_AGEMA_signal_3731 & n3915;
  LPM_q_ivl_22215 <= tmp_ivl_22217 & tmp_ivl_22212;
  new_AGEMA_signal_4041 <= tmp_ivl_22219(1);
  n3743 <= tmp_ivl_22219(0);
  tmp_ivl_22219 <= LPM_d0_ivl_22223(0 + 1 downto 0);
  tmp_ivl_22224 <= new_AGEMA_signal_4041 & n3743;
  LPM_q_ivl_22227 <= tmp_ivl_22229 & tmp_ivl_22224;
  tmp_ivl_22231 <= new_AGEMA_signal_4340 & n3742;
  LPM_q_ivl_22234 <= tmp_ivl_22236 & tmp_ivl_22231;
  tmp_ivl_22238 <= tmp_ivl_22242(1);
  tmp_ivl_22240 <= tmp_ivl_22242(0);
  tmp_ivl_22242 <= LPM_d0_ivl_22246(0 + 1 downto 0);
  tmp_ivl_22247 <= new_AGEMA_signal_3933 & n3745;
  LPM_q_ivl_22250 <= tmp_ivl_22252 & tmp_ivl_22247;
  tmp_ivl_22254 <= new_AGEMA_signal_3956 & n3744;
  LPM_q_ivl_22257 <= tmp_ivl_22259 & tmp_ivl_22254;
  new_AGEMA_signal_4341 <= tmp_ivl_22261(1);
  n3749 <= tmp_ivl_22261(0);
  tmp_ivl_22261 <= LPM_d0_ivl_22265(0 + 1 downto 0);
  tmp_ivl_22267 <= z1(5);
  tmp_ivl_22268 <= new_AGEMA_signal_3888 & tmp_ivl_22267;
  LPM_q_ivl_22271 <= tmp_ivl_22273 & tmp_ivl_22268;
  tmp_ivl_22276 <= state_in_s1(317);
  tmp_ivl_22278 <= state_in_s0(317);
  tmp_ivl_22279 <= tmp_ivl_22276 & tmp_ivl_22278;
  LPM_q_ivl_22282 <= tmp_ivl_22284 & tmp_ivl_22279;
  new_AGEMA_signal_4042 <= tmp_ivl_22286(1);
  n3748 <= tmp_ivl_22286(0);
  tmp_ivl_22286 <= LPM_d0_ivl_22290(0 + 1 downto 0);
  tmp_ivl_22292 <= state_in_s1(125);
  tmp_ivl_22294 <= state_in_s0(125);
  tmp_ivl_22295 <= tmp_ivl_22292 & tmp_ivl_22294;
  LPM_q_ivl_22298 <= tmp_ivl_22300 & tmp_ivl_22295;
  tmp_ivl_22302 <= new_AGEMA_signal_4039 & n3746;
  LPM_q_ivl_22305 <= tmp_ivl_22307 & tmp_ivl_22302;
  new_AGEMA_signal_4342 <= tmp_ivl_22309(1);
  n3747 <= tmp_ivl_22309(0);
  tmp_ivl_22309 <= LPM_d0_ivl_22313(0 + 1 downto 0);
  tmp_ivl_22314 <= new_AGEMA_signal_4042 & n3748;
  LPM_q_ivl_22317 <= tmp_ivl_22319 & tmp_ivl_22314;
  tmp_ivl_22321 <= new_AGEMA_signal_4342 & n3747;
  LPM_q_ivl_22324 <= tmp_ivl_22326 & tmp_ivl_22321;
  new_AGEMA_signal_4504 <= tmp_ivl_22328(1);
  n3755 <= tmp_ivl_22328(0);
  tmp_ivl_22328 <= LPM_d0_ivl_22332(0 + 1 downto 0);
  tmp_ivl_22333 <= new_AGEMA_signal_4341 & n3749;
  LPM_q_ivl_22336 <= tmp_ivl_22338 & tmp_ivl_22333;
  tmp_ivl_22340 <= new_AGEMA_signal_4504 & n3755;
  LPM_q_ivl_22343 <= tmp_ivl_22345 & tmp_ivl_22340;
  tmp_ivl_22347 <= tmp_ivl_22351(1);
  tmp_ivl_22349 <= tmp_ivl_22351(0);
  tmp_ivl_22351 <= LPM_d0_ivl_22355(0 + 1 downto 0);
  tmp_ivl_22356 <= new_AGEMA_signal_3932 & n3751;
  LPM_q_ivl_22359 <= tmp_ivl_22361 & tmp_ivl_22356;
  tmp_ivl_22363 <= new_AGEMA_signal_3935 & n3750;
  LPM_q_ivl_22366 <= tmp_ivl_22368 & tmp_ivl_22363;
  new_AGEMA_signal_4343 <= tmp_ivl_22370(1);
  n3752 <= tmp_ivl_22370(0);
  tmp_ivl_22370 <= LPM_d0_ivl_22374(0 + 1 downto 0);
  tmp_ivl_22375 <= new_AGEMA_signal_4343 & n3752;
  LPM_q_ivl_22378 <= tmp_ivl_22380 & tmp_ivl_22375;
  tmp_ivl_22382 <= new_AGEMA_signal_4504 & n3755;
  LPM_q_ivl_22385 <= tmp_ivl_22387 & tmp_ivl_22382;
  tmp_ivl_22389 <= tmp_ivl_22393(1);
  tmp_ivl_22391 <= tmp_ivl_22393(0);
  tmp_ivl_22393 <= LPM_d0_ivl_22397(0 + 1 downto 0);
  tmp_ivl_22398 <= new_AGEMA_signal_4029 & n3754;
  LPM_q_ivl_22401 <= tmp_ivl_22403 & tmp_ivl_22398;
  tmp_ivl_22405 <= new_AGEMA_signal_4586 & n3753;
  LPM_q_ivl_22408 <= tmp_ivl_22410 & tmp_ivl_22405;
  new_AGEMA_signal_4614 <= tmp_ivl_22412(1);
  n3756 <= tmp_ivl_22412(0);
  tmp_ivl_22412 <= LPM_d0_ivl_22416(0 + 1 downto 0);
  tmp_ivl_22417 <= new_AGEMA_signal_4614 & n3756;
  LPM_q_ivl_22420 <= tmp_ivl_22422 & tmp_ivl_22417;
  tmp_ivl_22424 <= new_AGEMA_signal_4504 & n3755;
  LPM_q_ivl_22427 <= tmp_ivl_22429 & tmp_ivl_22424;
  tmp_ivl_22431 <= tmp_ivl_22435(1);
  tmp_ivl_22433 <= tmp_ivl_22435(0);
  tmp_ivl_22435 <= LPM_d0_ivl_22439(0 + 1 downto 0);
  tmp_ivl_22440 <= new_AGEMA_signal_3732 & n3828;
  LPM_q_ivl_22443 <= tmp_ivl_22445 & tmp_ivl_22440;
  tmp_ivl_22447 <= new_AGEMA_signal_3742 & n3914;
  LPM_q_ivl_22450 <= tmp_ivl_22452 & tmp_ivl_22447;
  new_AGEMA_signal_4043 <= tmp_ivl_22454(1);
  n3758 <= tmp_ivl_22454(0);
  tmp_ivl_22454 <= LPM_d0_ivl_22458(0 + 1 downto 0);
  tmp_ivl_22460 <= z0(6);
  tmp_ivl_22461 <= new_AGEMA_signal_4202 & tmp_ivl_22460;
  LPM_q_ivl_22464 <= tmp_ivl_22466 & tmp_ivl_22461;
  tmp_ivl_22469 <= state_in_s1(62);
  tmp_ivl_22471 <= state_in_s0(62);
  tmp_ivl_22472 <= tmp_ivl_22469 & tmp_ivl_22471;
  LPM_q_ivl_22475 <= tmp_ivl_22477 & tmp_ivl_22472;
  new_AGEMA_signal_4344 <= tmp_ivl_22479(1);
  n3763 <= tmp_ivl_22479(0);
  tmp_ivl_22479 <= LPM_d0_ivl_22483(0 + 1 downto 0);
  tmp_ivl_22484 <= new_AGEMA_signal_4344 & n3763;
  LPM_q_ivl_22487 <= tmp_ivl_22489 & tmp_ivl_22484;
  tmp_ivl_22491 <= new_AGEMA_signal_3319 & n3757;
  LPM_q_ivl_22494 <= tmp_ivl_22496 & tmp_ivl_22491;
  new_AGEMA_signal_4505 <= tmp_ivl_22498(1);
  n3822 <= tmp_ivl_22498(0);
  tmp_ivl_22498 <= LPM_d0_ivl_22502(0 + 1 downto 0);
  tmp_ivl_22503 <= new_AGEMA_signal_4043 & n3758;
  LPM_q_ivl_22506 <= tmp_ivl_22508 & tmp_ivl_22503;
  tmp_ivl_22510 <= new_AGEMA_signal_4505 & n3822;
  LPM_q_ivl_22513 <= tmp_ivl_22515 & tmp_ivl_22510;
  tmp_ivl_22517 <= tmp_ivl_22521(1);
  tmp_ivl_22519 <= tmp_ivl_22521(0);
  tmp_ivl_22521 <= LPM_d0_ivl_22525(0 + 1 downto 0);
  tmp_ivl_22526 <= new_AGEMA_signal_3716 & n3760;
  LPM_q_ivl_22529 <= tmp_ivl_22531 & tmp_ivl_22526;
  tmp_ivl_22533 <= new_AGEMA_signal_3744 & n3759;
  LPM_q_ivl_22536 <= tmp_ivl_22538 & tmp_ivl_22533;
  new_AGEMA_signal_4044 <= tmp_ivl_22540(1);
  n3761 <= tmp_ivl_22540(0);
  tmp_ivl_22540 <= LPM_d0_ivl_22544(0 + 1 downto 0);
  tmp_ivl_22545 <= new_AGEMA_signal_4044 & n3761;
  LPM_q_ivl_22548 <= tmp_ivl_22550 & tmp_ivl_22545;
  tmp_ivl_22552 <= new_AGEMA_signal_4505 & n3822;
  LPM_q_ivl_22555 <= tmp_ivl_22557 & tmp_ivl_22552;
  tmp_ivl_22559 <= tmp_ivl_22563(1);
  tmp_ivl_22561 <= tmp_ivl_22563(0);
  tmp_ivl_22563 <= LPM_d0_ivl_22567(0 + 1 downto 0);
  tmp_ivl_22568 <= new_AGEMA_signal_3941 & n3762;
  LPM_q_ivl_22571 <= tmp_ivl_22573 & tmp_ivl_22568;
  tmp_ivl_22575 <= new_AGEMA_signal_3966 & n3809;
  LPM_q_ivl_22578 <= tmp_ivl_22580 & tmp_ivl_22575;
  new_AGEMA_signal_4345 <= tmp_ivl_22582(1);
  n3766 <= tmp_ivl_22582(0);
  tmp_ivl_22582 <= LPM_d0_ivl_22586(0 + 1 downto 0);
  tmp_ivl_22588 <= z1(6);
  tmp_ivl_22589 <= new_AGEMA_signal_4201 & tmp_ivl_22588;
  LPM_q_ivl_22592 <= tmp_ivl_22594 & tmp_ivl_22589;
  tmp_ivl_22597 <= state_in_s1(318);
  tmp_ivl_22599 <= state_in_s0(318);
  tmp_ivl_22600 <= tmp_ivl_22597 & tmp_ivl_22599;
  LPM_q_ivl_22603 <= tmp_ivl_22605 & tmp_ivl_22600;
  new_AGEMA_signal_4346 <= tmp_ivl_22607(1);
  n3765 <= tmp_ivl_22607(0);
  tmp_ivl_22607 <= LPM_d0_ivl_22611(0 + 1 downto 0);
  tmp_ivl_22613 <= state_in_s1(126);
  tmp_ivl_22615 <= state_in_s0(126);
  tmp_ivl_22616 <= tmp_ivl_22613 & tmp_ivl_22615;
  LPM_q_ivl_22619 <= tmp_ivl_22621 & tmp_ivl_22616;
  tmp_ivl_22623 <= new_AGEMA_signal_4344 & n3763;
  LPM_q_ivl_22626 <= tmp_ivl_22628 & tmp_ivl_22623;
  new_AGEMA_signal_4506 <= tmp_ivl_22630(1);
  n3764 <= tmp_ivl_22630(0);
  tmp_ivl_22630 <= LPM_d0_ivl_22634(0 + 1 downto 0);
  tmp_ivl_22635 <= new_AGEMA_signal_4346 & n3765;
  LPM_q_ivl_22638 <= tmp_ivl_22640 & tmp_ivl_22635;
  tmp_ivl_22642 <= new_AGEMA_signal_4506 & n3764;
  LPM_q_ivl_22645 <= tmp_ivl_22647 & tmp_ivl_22642;
  new_AGEMA_signal_4591 <= tmp_ivl_22649(1);
  n3819 <= tmp_ivl_22649(0);
  tmp_ivl_22649 <= LPM_d0_ivl_22653(0 + 1 downto 0);
  tmp_ivl_22654 <= new_AGEMA_signal_4345 & n3766;
  LPM_q_ivl_22657 <= tmp_ivl_22659 & tmp_ivl_22654;
  tmp_ivl_22661 <= new_AGEMA_signal_4591 & n3819;
  LPM_q_ivl_22664 <= tmp_ivl_22666 & tmp_ivl_22661;
  tmp_ivl_22668 <= tmp_ivl_22672(1);
  tmp_ivl_22670 <= tmp_ivl_22672(0);
  tmp_ivl_22672 <= LPM_d0_ivl_22676(0 + 1 downto 0);
  tmp_ivl_22677 <= new_AGEMA_signal_3940 & n3767;
  LPM_q_ivl_22680 <= tmp_ivl_22682 & tmp_ivl_22677;
  tmp_ivl_22684 <= new_AGEMA_signal_3943 & n3791;
  LPM_q_ivl_22687 <= tmp_ivl_22689 & tmp_ivl_22684;
  new_AGEMA_signal_4347 <= tmp_ivl_22691(1);
  n3768 <= tmp_ivl_22691(0);
  tmp_ivl_22691 <= LPM_d0_ivl_22695(0 + 1 downto 0);
  tmp_ivl_22696 <= new_AGEMA_signal_4347 & n3768;
  LPM_q_ivl_22699 <= tmp_ivl_22701 & tmp_ivl_22696;
  tmp_ivl_22703 <= new_AGEMA_signal_4591 & n3819;
  LPM_q_ivl_22706 <= tmp_ivl_22708 & tmp_ivl_22703;
  tmp_ivl_22710 <= tmp_ivl_22714(1);
  tmp_ivl_22712 <= tmp_ivl_22714(0);
  tmp_ivl_22714 <= LPM_d0_ivl_22718(0 + 1 downto 0);
  tmp_ivl_22719 <= new_AGEMA_signal_3382 & n3770;
  LPM_q_ivl_22722 <= tmp_ivl_22724 & tmp_ivl_22719;
  tmp_ivl_22726 <= new_AGEMA_signal_3375 & n3769;
  LPM_q_ivl_22729 <= tmp_ivl_22731 & tmp_ivl_22726;
  new_AGEMA_signal_3750 <= tmp_ivl_22733(1);
  n3875 <= tmp_ivl_22733(0);
  tmp_ivl_22733 <= LPM_d0_ivl_22737(0 + 1 downto 0);
  tmp_ivl_22738 <= new_AGEMA_signal_3714 & n3872;
  LPM_q_ivl_22741 <= tmp_ivl_22743 & tmp_ivl_22738;
  tmp_ivl_22745 <= new_AGEMA_signal_3750 & n3875;
  LPM_q_ivl_22748 <= tmp_ivl_22750 & tmp_ivl_22745;
  new_AGEMA_signal_4045 <= tmp_ivl_22752(1);
  n3772 <= tmp_ivl_22752(0);
  tmp_ivl_22752 <= LPM_d0_ivl_22756(0 + 1 downto 0);
  tmp_ivl_22758 <= state_in_s1(233);
  tmp_ivl_22760 <= state_in_s0(233);
  tmp_ivl_22761 <= tmp_ivl_22758 & tmp_ivl_22760;
  LPM_q_ivl_22764 <= tmp_ivl_22766 & tmp_ivl_22761;
  tmp_ivl_22769 <= z4(17);
  tmp_ivl_22770 <= new_AGEMA_signal_3119 & tmp_ivl_22769;
  LPM_q_ivl_22773 <= tmp_ivl_22775 & tmp_ivl_22770;
  new_AGEMA_signal_3447 <= tmp_ivl_22777(1);
  n3778 <= tmp_ivl_22777(0);
  tmp_ivl_22777 <= LPM_d0_ivl_22781(0 + 1 downto 0);
  tmp_ivl_22782 <= new_AGEMA_signal_3361 & n3771;
  LPM_q_ivl_22785 <= tmp_ivl_22787 & tmp_ivl_22782;
  tmp_ivl_22789 <= new_AGEMA_signal_3447 & n3778;
  LPM_q_ivl_22792 <= tmp_ivl_22794 & tmp_ivl_22789;
  new_AGEMA_signal_3751 <= tmp_ivl_22796(1);
  n3786 <= tmp_ivl_22796(0);
  tmp_ivl_22796 <= LPM_d0_ivl_22800(0 + 1 downto 0);
  tmp_ivl_22801 <= new_AGEMA_signal_4045 & n3772;
  LPM_q_ivl_22804 <= tmp_ivl_22806 & tmp_ivl_22801;
  tmp_ivl_22808 <= new_AGEMA_signal_3751 & n3786;
  LPM_q_ivl_22811 <= tmp_ivl_22813 & tmp_ivl_22808;
  tmp_ivl_22815 <= tmp_ivl_22819(1);
  tmp_ivl_22817 <= tmp_ivl_22819(0);
  tmp_ivl_22819 <= LPM_d0_ivl_22823(0 + 1 downto 0);
  tmp_ivl_22824 <= new_AGEMA_signal_3673 & n3774;
  LPM_q_ivl_22827 <= tmp_ivl_22829 & tmp_ivl_22824;
  tmp_ivl_22831 <= new_AGEMA_signal_3715 & n3773;
  LPM_q_ivl_22834 <= tmp_ivl_22836 & tmp_ivl_22831;
  new_AGEMA_signal_4046 <= tmp_ivl_22838(1);
  n3775 <= tmp_ivl_22838(0);
  tmp_ivl_22838 <= LPM_d0_ivl_22842(0 + 1 downto 0);
  tmp_ivl_22843 <= new_AGEMA_signal_4046 & n3775;
  LPM_q_ivl_22846 <= tmp_ivl_22848 & tmp_ivl_22843;
  tmp_ivl_22850 <= new_AGEMA_signal_3751 & n3786;
  LPM_q_ivl_22853 <= tmp_ivl_22855 & tmp_ivl_22850;
  tmp_ivl_22857 <= tmp_ivl_22861(1);
  tmp_ivl_22859 <= tmp_ivl_22861(0);
  tmp_ivl_22861 <= LPM_d0_ivl_22865(0 + 1 downto 0);
  tmp_ivl_22866 <= new_AGEMA_signal_3608 & n3777;
  LPM_q_ivl_22869 <= tmp_ivl_22871 & tmp_ivl_22866;
  tmp_ivl_22873 <= new_AGEMA_signal_3612 & n3776;
  LPM_q_ivl_22876 <= tmp_ivl_22878 & tmp_ivl_22873;
  new_AGEMA_signal_4047 <= tmp_ivl_22880(1);
  n3779 <= tmp_ivl_22880(0);
  tmp_ivl_22880 <= LPM_d0_ivl_22884(0 + 1 downto 0);
  tmp_ivl_22886 <= state_in_s1(297);
  tmp_ivl_22888 <= state_in_s0(297);
  tmp_ivl_22889 <= tmp_ivl_22886 & tmp_ivl_22888;
  LPM_q_ivl_22892 <= tmp_ivl_22894 & tmp_ivl_22889;
  tmp_ivl_22896 <= new_AGEMA_signal_3447 & n3778;
  LPM_q_ivl_22899 <= tmp_ivl_22901 & tmp_ivl_22896;
  new_AGEMA_signal_3752 <= tmp_ivl_22903(1);
  n3838 <= tmp_ivl_22903(0);
  tmp_ivl_22903 <= LPM_d0_ivl_22907(0 + 1 downto 0);
  tmp_ivl_22908 <= new_AGEMA_signal_4047 & n3779;
  LPM_q_ivl_22911 <= tmp_ivl_22913 & tmp_ivl_22908;
  tmp_ivl_22915 <= new_AGEMA_signal_3752 & n3838;
  LPM_q_ivl_22918 <= tmp_ivl_22920 & tmp_ivl_22915;
  tmp_ivl_22922 <= tmp_ivl_22926(1);
  tmp_ivl_22924 <= tmp_ivl_22926(0);
  tmp_ivl_22926 <= LPM_d0_ivl_22930(0 + 1 downto 0);
  tmp_ivl_22931 <= new_AGEMA_signal_3639 & n3780;
  LPM_q_ivl_22934 <= tmp_ivl_22936 & tmp_ivl_22931;
  tmp_ivl_22938 <= new_AGEMA_signal_3642 & n3832;
  LPM_q_ivl_22941 <= tmp_ivl_22943 & tmp_ivl_22938;
  new_AGEMA_signal_4048 <= tmp_ivl_22945(1);
  n3781 <= tmp_ivl_22945(0);
  tmp_ivl_22945 <= LPM_d0_ivl_22949(0 + 1 downto 0);
  tmp_ivl_22950 <= new_AGEMA_signal_4048 & n3781;
  LPM_q_ivl_22953 <= tmp_ivl_22955 & tmp_ivl_22950;
  tmp_ivl_22957 <= new_AGEMA_signal_3752 & n3838;
  LPM_q_ivl_22960 <= tmp_ivl_22962 & tmp_ivl_22957;
  tmp_ivl_22964 <= tmp_ivl_22968(1);
  tmp_ivl_22966 <= tmp_ivl_22968(0);
  tmp_ivl_22968 <= LPM_d0_ivl_22972(0 + 1 downto 0);
  tmp_ivl_22973 <= new_AGEMA_signal_3689 & n3860;
  LPM_q_ivl_22976 <= tmp_ivl_22978 & tmp_ivl_22973;
  tmp_ivl_22980 <= new_AGEMA_signal_4009 & n3782;
  LPM_q_ivl_22983 <= tmp_ivl_22985 & tmp_ivl_22980;
  new_AGEMA_signal_4352 <= tmp_ivl_22987(1);
  n3784 <= tmp_ivl_22987(0);
  tmp_ivl_22987 <= LPM_d0_ivl_22991(0 + 1 downto 0);
  tmp_ivl_22993 <= z0(45);
  tmp_ivl_22994 <= new_AGEMA_signal_3214 & tmp_ivl_22993;
  LPM_q_ivl_22997 <= tmp_ivl_22999 & tmp_ivl_22994;
  tmp_ivl_23002 <= state_in_s1(21);
  tmp_ivl_23004 <= state_in_s0(21);
  tmp_ivl_23005 <= tmp_ivl_23002 & tmp_ivl_23004;
  LPM_q_ivl_23008 <= tmp_ivl_23010 & tmp_ivl_23005;
  new_AGEMA_signal_3448 <= tmp_ivl_23012(1);
  n3792 <= tmp_ivl_23012(0);
  tmp_ivl_23012 <= LPM_d0_ivl_23016(0 + 1 downto 0);
  tmp_ivl_23017 <= new_AGEMA_signal_3448 & n3792;
  LPM_q_ivl_23020 <= tmp_ivl_23022 & tmp_ivl_23017;
  tmp_ivl_23024 <= new_AGEMA_signal_3308 & n3783;
  LPM_q_ivl_23027 <= tmp_ivl_23029 & tmp_ivl_23024;
  new_AGEMA_signal_3753 <= tmp_ivl_23031(1);
  n3788 <= tmp_ivl_23031(0);
  tmp_ivl_23031 <= LPM_d0_ivl_23035(0 + 1 downto 0);
  tmp_ivl_23036 <= new_AGEMA_signal_4352 & n3784;
  LPM_q_ivl_23039 <= tmp_ivl_23041 & tmp_ivl_23036;
  tmp_ivl_23043 <= new_AGEMA_signal_3753 & n3788;
  LPM_q_ivl_23046 <= tmp_ivl_23048 & tmp_ivl_23043;
  tmp_ivl_23050 <= tmp_ivl_23054(1);
  tmp_ivl_23052 <= tmp_ivl_23054(0);
  tmp_ivl_23054 <= LPM_d0_ivl_23058(0 + 1 downto 0);
  tmp_ivl_23059 <= new_AGEMA_signal_3720 & n3859;
  LPM_q_ivl_23062 <= tmp_ivl_23064 & tmp_ivl_23059;
  tmp_ivl_23066 <= new_AGEMA_signal_3750 & n3875;
  LPM_q_ivl_23069 <= tmp_ivl_23071 & tmp_ivl_23066;
  new_AGEMA_signal_4049 <= tmp_ivl_23073(1);
  n3785 <= tmp_ivl_23073(0);
  tmp_ivl_23073 <= LPM_d0_ivl_23077(0 + 1 downto 0);
  tmp_ivl_23078 <= new_AGEMA_signal_4049 & n3785;
  LPM_q_ivl_23081 <= tmp_ivl_23083 & tmp_ivl_23078;
  tmp_ivl_23085 <= new_AGEMA_signal_3753 & n3788;
  LPM_q_ivl_23088 <= tmp_ivl_23090 & tmp_ivl_23085;
  tmp_ivl_23092 <= tmp_ivl_23096(1);
  tmp_ivl_23094 <= tmp_ivl_23096(0);
  tmp_ivl_23096 <= LPM_d0_ivl_23100(0 + 1 downto 0);
  tmp_ivl_23101 <= new_AGEMA_signal_3672 & n3787;
  LPM_q_ivl_23104 <= tmp_ivl_23106 & tmp_ivl_23101;
  tmp_ivl_23108 <= new_AGEMA_signal_3751 & n3786;
  LPM_q_ivl_23111 <= tmp_ivl_23113 & tmp_ivl_23108;
  new_AGEMA_signal_4050 <= tmp_ivl_23115(1);
  n3789 <= tmp_ivl_23115(0);
  tmp_ivl_23115 <= LPM_d0_ivl_23119(0 + 1 downto 0);
  tmp_ivl_23120 <= new_AGEMA_signal_4050 & n3789;
  LPM_q_ivl_23123 <= tmp_ivl_23125 & tmp_ivl_23120;
  tmp_ivl_23127 <= new_AGEMA_signal_3753 & n3788;
  LPM_q_ivl_23130 <= tmp_ivl_23132 & tmp_ivl_23127;
  tmp_ivl_23134 <= tmp_ivl_23138(1);
  tmp_ivl_23136 <= tmp_ivl_23138(0);
  tmp_ivl_23138 <= LPM_d0_ivl_23142(0 + 1 downto 0);
  tmp_ivl_23143 <= new_AGEMA_signal_3943 & n3791;
  LPM_q_ivl_23146 <= tmp_ivl_23148 & tmp_ivl_23143;
  tmp_ivl_23150 <= new_AGEMA_signal_3994 & n3790;
  LPM_q_ivl_23153 <= tmp_ivl_23155 & tmp_ivl_23150;
  new_AGEMA_signal_4355 <= tmp_ivl_23157(1);
  n3795 <= tmp_ivl_23157(0);
  tmp_ivl_23157 <= LPM_d0_ivl_23161(0 + 1 downto 0);
  tmp_ivl_23163 <= z1(45);
  tmp_ivl_23164 <= new_AGEMA_signal_3026 & tmp_ivl_23163;
  LPM_q_ivl_23167 <= tmp_ivl_23169 & tmp_ivl_23164;
  tmp_ivl_23171 <= new_AGEMA_signal_3448 & n3792;
  LPM_q_ivl_23174 <= tmp_ivl_23176 & tmp_ivl_23171;
  new_AGEMA_signal_3754 <= tmp_ivl_23178(1);
  n3794 <= tmp_ivl_23178(0);
  tmp_ivl_23178 <= LPM_d0_ivl_23182(0 + 1 downto 0);
  tmp_ivl_23183 <= new_AGEMA_signal_3754 & n3794;
  LPM_q_ivl_23186 <= tmp_ivl_23188 & tmp_ivl_23183;
  tmp_ivl_23190 <= new_AGEMA_signal_2689 & n3793;
  LPM_q_ivl_23193 <= tmp_ivl_23195 & tmp_ivl_23190;
  new_AGEMA_signal_4051 <= tmp_ivl_23197(1);
  n3818 <= tmp_ivl_23197(0);
  tmp_ivl_23197 <= LPM_d0_ivl_23201(0 + 1 downto 0);
  tmp_ivl_23202 <= new_AGEMA_signal_4355 & n3795;
  LPM_q_ivl_23205 <= tmp_ivl_23207 & tmp_ivl_23202;
  tmp_ivl_23209 <= new_AGEMA_signal_4051 & n3818;
  LPM_q_ivl_23212 <= tmp_ivl_23214 & tmp_ivl_23209;
  tmp_ivl_23216 <= tmp_ivl_23220(1);
  tmp_ivl_23218 <= tmp_ivl_23220(0);
  tmp_ivl_23220 <= LPM_d0_ivl_23224(0 + 1 downto 0);
  tmp_ivl_23225 <= new_AGEMA_signal_3925 & n3796;
  LPM_q_ivl_23228 <= tmp_ivl_23230 & tmp_ivl_23225;
  tmp_ivl_23232 <= new_AGEMA_signal_4003 & n3816;
  LPM_q_ivl_23235 <= tmp_ivl_23237 & tmp_ivl_23232;
  new_AGEMA_signal_4356 <= tmp_ivl_23239(1);
  n3797 <= tmp_ivl_23239(0);
  tmp_ivl_23239 <= LPM_d0_ivl_23243(0 + 1 downto 0);
  tmp_ivl_23244 <= new_AGEMA_signal_4356 & n3797;
  LPM_q_ivl_23247 <= tmp_ivl_23249 & tmp_ivl_23244;
  tmp_ivl_23251 <= new_AGEMA_signal_4051 & n3818;
  LPM_q_ivl_23254 <= tmp_ivl_23256 & tmp_ivl_23251;
  tmp_ivl_23258 <= tmp_ivl_23262(1);
  tmp_ivl_23260 <= tmp_ivl_23262(0);
  tmp_ivl_23262 <= LPM_d0_ivl_23266(0 + 1 downto 0);
  tmp_ivl_23267 <= new_AGEMA_signal_3695 & n3799;
  LPM_q_ivl_23270 <= tmp_ivl_23272 & tmp_ivl_23267;
  tmp_ivl_23274 <= new_AGEMA_signal_3704 & n3798;
  LPM_q_ivl_23277 <= tmp_ivl_23279 & tmp_ivl_23274;
  new_AGEMA_signal_4052 <= tmp_ivl_23281(1);
  n3801 <= tmp_ivl_23281(0);
  tmp_ivl_23281 <= LPM_d0_ivl_23285(0 + 1 downto 0);
  tmp_ivl_23287 <= z0(3);
  tmp_ivl_23288 <= new_AGEMA_signal_4580 & tmp_ivl_23287;
  LPM_q_ivl_23291 <= tmp_ivl_23293 & tmp_ivl_23288;
  tmp_ivl_23296 <= state_in_s1(59);
  tmp_ivl_23298 <= state_in_s0(59);
  tmp_ivl_23299 <= tmp_ivl_23296 & tmp_ivl_23298;
  LPM_q_ivl_23302 <= tmp_ivl_23304 & tmp_ivl_23299;
  new_AGEMA_signal_4592 <= tmp_ivl_23306(1);
  n3811 <= tmp_ivl_23306(0);
  tmp_ivl_23306 <= LPM_d0_ivl_23310(0 + 1 downto 0);
  tmp_ivl_23311 <= new_AGEMA_signal_4592 & n3811;
  LPM_q_ivl_23314 <= tmp_ivl_23316 & tmp_ivl_23311;
  tmp_ivl_23318 <= new_AGEMA_signal_3306 & n3800;
  LPM_q_ivl_23321 <= tmp_ivl_23323 & tmp_ivl_23318;
  new_AGEMA_signal_4617 <= tmp_ivl_23325(1);
  n3807 <= tmp_ivl_23325(0);
  tmp_ivl_23325 <= LPM_d0_ivl_23329(0 + 1 downto 0);
  tmp_ivl_23330 <= new_AGEMA_signal_4052 & n3801;
  LPM_q_ivl_23333 <= tmp_ivl_23335 & tmp_ivl_23330;
  tmp_ivl_23337 <= new_AGEMA_signal_4617 & n3807;
  LPM_q_ivl_23340 <= tmp_ivl_23342 & tmp_ivl_23337;
  tmp_ivl_23344 <= tmp_ivl_23348(1);
  tmp_ivl_23346 <= tmp_ivl_23348(0);
  tmp_ivl_23348 <= LPM_d0_ivl_23352(0 + 1 downto 0);
  tmp_ivl_23353 <= new_AGEMA_signal_3668 & n3803;
  LPM_q_ivl_23356 <= tmp_ivl_23358 & tmp_ivl_23353;
  tmp_ivl_23360 <= new_AGEMA_signal_3703 & n3802;
  LPM_q_ivl_23363 <= tmp_ivl_23365 & tmp_ivl_23360;
  new_AGEMA_signal_4053 <= tmp_ivl_23367(1);
  n3804 <= tmp_ivl_23367(0);
  tmp_ivl_23367 <= LPM_d0_ivl_23371(0 + 1 downto 0);
  tmp_ivl_23372 <= new_AGEMA_signal_4053 & n3804;
  LPM_q_ivl_23375 <= tmp_ivl_23377 & tmp_ivl_23372;
  tmp_ivl_23379 <= new_AGEMA_signal_4617 & n3807;
  LPM_q_ivl_23382 <= tmp_ivl_23384 & tmp_ivl_23379;
  tmp_ivl_23386 <= tmp_ivl_23390(1);
  tmp_ivl_23388 <= tmp_ivl_23390(0);
  tmp_ivl_23390 <= LPM_d0_ivl_23394(0 + 1 downto 0);
  tmp_ivl_23395 <= new_AGEMA_signal_3667 & n3806;
  LPM_q_ivl_23398 <= tmp_ivl_23400 & tmp_ivl_23395;
  tmp_ivl_23402 <= new_AGEMA_signal_3711 & n3805;
  LPM_q_ivl_23405 <= tmp_ivl_23407 & tmp_ivl_23402;
  new_AGEMA_signal_4054 <= tmp_ivl_23409(1);
  n3808 <= tmp_ivl_23409(0);
  tmp_ivl_23409 <= LPM_d0_ivl_23413(0 + 1 downto 0);
  tmp_ivl_23414 <= new_AGEMA_signal_4054 & n3808;
  LPM_q_ivl_23417 <= tmp_ivl_23419 & tmp_ivl_23414;
  tmp_ivl_23421 <= new_AGEMA_signal_4617 & n3807;
  LPM_q_ivl_23424 <= tmp_ivl_23426 & tmp_ivl_23421;
  tmp_ivl_23428 <= tmp_ivl_23432(1);
  tmp_ivl_23430 <= tmp_ivl_23432(0);
  tmp_ivl_23432 <= LPM_d0_ivl_23436(0 + 1 downto 0);
  tmp_ivl_23437 <= new_AGEMA_signal_3934 & n3810;
  LPM_q_ivl_23440 <= tmp_ivl_23442 & tmp_ivl_23437;
  tmp_ivl_23444 <= new_AGEMA_signal_3966 & n3809;
  LPM_q_ivl_23447 <= tmp_ivl_23449 & tmp_ivl_23444;
  new_AGEMA_signal_4357 <= tmp_ivl_23451(1);
  n3814 <= tmp_ivl_23451(0);
  tmp_ivl_23451 <= LPM_d0_ivl_23455(0 + 1 downto 0);
  tmp_ivl_23457 <= z1(3);
  tmp_ivl_23458 <= new_AGEMA_signal_4577 & tmp_ivl_23457;
  LPM_q_ivl_23461 <= tmp_ivl_23463 & tmp_ivl_23458;
  tmp_ivl_23466 <= state_in_s1(315);
  tmp_ivl_23468 <= state_in_s0(315);
  tmp_ivl_23469 <= tmp_ivl_23466 & tmp_ivl_23468;
  LPM_q_ivl_23472 <= tmp_ivl_23474 & tmp_ivl_23469;
  new_AGEMA_signal_4593 <= tmp_ivl_23476(1);
  n3813 <= tmp_ivl_23476(0);
  tmp_ivl_23476 <= LPM_d0_ivl_23480(0 + 1 downto 0);
  tmp_ivl_23482 <= state_in_s1(123);
  tmp_ivl_23484 <= state_in_s0(123);
  tmp_ivl_23485 <= tmp_ivl_23482 & tmp_ivl_23484;
  LPM_q_ivl_23488 <= tmp_ivl_23490 & tmp_ivl_23485;
  tmp_ivl_23492 <= new_AGEMA_signal_4592 & n3811;
  LPM_q_ivl_23495 <= tmp_ivl_23497 & tmp_ivl_23492;
  new_AGEMA_signal_4618 <= tmp_ivl_23499(1);
  n3812 <= tmp_ivl_23499(0);
  tmp_ivl_23499 <= LPM_d0_ivl_23503(0 + 1 downto 0);
  tmp_ivl_23504 <= new_AGEMA_signal_4593 & n3813;
  LPM_q_ivl_23507 <= tmp_ivl_23509 & tmp_ivl_23504;
  tmp_ivl_23511 <= new_AGEMA_signal_4618 & n3812;
  LPM_q_ivl_23514 <= tmp_ivl_23516 & tmp_ivl_23511;
  new_AGEMA_signal_4639 <= tmp_ivl_23518(1);
  n3820 <= tmp_ivl_23518(0);
  tmp_ivl_23518 <= LPM_d0_ivl_23522(0 + 1 downto 0);
  tmp_ivl_23523 <= new_AGEMA_signal_4357 & n3814;
  LPM_q_ivl_23526 <= tmp_ivl_23528 & tmp_ivl_23523;
  tmp_ivl_23530 <= new_AGEMA_signal_4639 & n3820;
  LPM_q_ivl_23533 <= tmp_ivl_23535 & tmp_ivl_23530;
  tmp_ivl_23537 <= tmp_ivl_23541(1);
  tmp_ivl_23539 <= tmp_ivl_23541(0);
  tmp_ivl_23541 <= LPM_d0_ivl_23545(0 + 1 downto 0);
  tmp_ivl_23546 <= new_AGEMA_signal_4003 & n3816;
  LPM_q_ivl_23549 <= tmp_ivl_23551 & tmp_ivl_23546;
  tmp_ivl_23553 <= new_AGEMA_signal_4310 & n3815;
  LPM_q_ivl_23556 <= tmp_ivl_23558 & tmp_ivl_23553;
  new_AGEMA_signal_4510 <= tmp_ivl_23560(1);
  n3817 <= tmp_ivl_23560(0);
  tmp_ivl_23560 <= LPM_d0_ivl_23564(0 + 1 downto 0);
  tmp_ivl_23565 <= new_AGEMA_signal_4510 & n3817;
  LPM_q_ivl_23568 <= tmp_ivl_23570 & tmp_ivl_23565;
  tmp_ivl_23572 <= new_AGEMA_signal_4639 & n3820;
  LPM_q_ivl_23575 <= tmp_ivl_23577 & tmp_ivl_23572;
  tmp_ivl_23579 <= tmp_ivl_23583(1);
  tmp_ivl_23581 <= tmp_ivl_23583(0);
  tmp_ivl_23583 <= LPM_d0_ivl_23587(0 + 1 downto 0);
  tmp_ivl_23588 <= new_AGEMA_signal_4591 & n3819;
  LPM_q_ivl_23591 <= tmp_ivl_23593 & tmp_ivl_23588;
  tmp_ivl_23595 <= new_AGEMA_signal_4051 & n3818;
  LPM_q_ivl_23598 <= tmp_ivl_23600 & tmp_ivl_23595;
  new_AGEMA_signal_4619 <= tmp_ivl_23602(1);
  n3821 <= tmp_ivl_23602(0);
  tmp_ivl_23602 <= LPM_d0_ivl_23606(0 + 1 downto 0);
  tmp_ivl_23607 <= new_AGEMA_signal_4619 & n3821;
  LPM_q_ivl_23610 <= tmp_ivl_23612 & tmp_ivl_23607;
  tmp_ivl_23614 <= new_AGEMA_signal_4639 & n3820;
  LPM_q_ivl_23617 <= tmp_ivl_23619 & tmp_ivl_23614;
  tmp_ivl_23621 <= tmp_ivl_23625(1);
  tmp_ivl_23623 <= tmp_ivl_23625(0);
  tmp_ivl_23625 <= LPM_d0_ivl_23629(0 + 1 downto 0);
  tmp_ivl_23630 <= new_AGEMA_signal_3693 & n3823;
  LPM_q_ivl_23633 <= tmp_ivl_23635 & tmp_ivl_23630;
  tmp_ivl_23637 <= new_AGEMA_signal_4505 & n3822;
  LPM_q_ivl_23640 <= tmp_ivl_23642 & tmp_ivl_23637;
  new_AGEMA_signal_4594 <= tmp_ivl_23644(1);
  n3825 <= tmp_ivl_23644(0);
  tmp_ivl_23644 <= LPM_d0_ivl_23648(0 + 1 downto 0);
  tmp_ivl_23650 <= state_in_s1(203);
  tmp_ivl_23652 <= state_in_s0(203);
  tmp_ivl_23653 <= tmp_ivl_23650 & tmp_ivl_23652;
  LPM_q_ivl_23656 <= tmp_ivl_23658 & tmp_ivl_23653;
  tmp_ivl_23661 <= z4(51);
  tmp_ivl_23662 <= new_AGEMA_signal_3157 & tmp_ivl_23661;
  LPM_q_ivl_23665 <= tmp_ivl_23667 & tmp_ivl_23662;
  new_AGEMA_signal_3449 <= tmp_ivl_23669(1);
  n3833 <= tmp_ivl_23669(0);
  tmp_ivl_23669 <= LPM_d0_ivl_23673(0 + 1 downto 0);
  tmp_ivl_23674 <= new_AGEMA_signal_3384 & n3824;
  LPM_q_ivl_23677 <= tmp_ivl_23679 & tmp_ivl_23674;
  tmp_ivl_23681 <= new_AGEMA_signal_3449 & n3833;
  LPM_q_ivl_23684 <= tmp_ivl_23686 & tmp_ivl_23681;
  new_AGEMA_signal_3755 <= tmp_ivl_23688(1);
  n3829 <= tmp_ivl_23688(0);
  tmp_ivl_23688 <= LPM_d0_ivl_23692(0 + 1 downto 0);
  tmp_ivl_23693 <= new_AGEMA_signal_4594 & n3825;
  LPM_q_ivl_23696 <= tmp_ivl_23698 & tmp_ivl_23693;
  tmp_ivl_23700 <= new_AGEMA_signal_3755 & n3829;
  LPM_q_ivl_23703 <= tmp_ivl_23705 & tmp_ivl_23700;
  tmp_ivl_23707 <= tmp_ivl_23711(1);
  tmp_ivl_23709 <= tmp_ivl_23711(0);
  tmp_ivl_23711 <= LPM_d0_ivl_23715(0 + 1 downto 0);
  tmp_ivl_23716 <= new_AGEMA_signal_3692 & n3826;
  LPM_q_ivl_23719 <= tmp_ivl_23721 & tmp_ivl_23716;
  tmp_ivl_23723 <= new_AGEMA_signal_3728 & n3893;
  LPM_q_ivl_23726 <= tmp_ivl_23728 & tmp_ivl_23723;
  new_AGEMA_signal_4055 <= tmp_ivl_23730(1);
  n3827 <= tmp_ivl_23730(0);
  tmp_ivl_23730 <= LPM_d0_ivl_23734(0 + 1 downto 0);
  tmp_ivl_23735 <= new_AGEMA_signal_4055 & n3827;
  LPM_q_ivl_23738 <= tmp_ivl_23740 & tmp_ivl_23735;
  tmp_ivl_23742 <= new_AGEMA_signal_3755 & n3829;
  LPM_q_ivl_23745 <= tmp_ivl_23747 & tmp_ivl_23742;
  tmp_ivl_23749 <= tmp_ivl_23753(1);
  tmp_ivl_23751 <= tmp_ivl_23753(0);
  tmp_ivl_23753 <= LPM_d0_ivl_23757(0 + 1 downto 0);
  tmp_ivl_23758 <= new_AGEMA_signal_3724 & n3894;
  LPM_q_ivl_23761 <= tmp_ivl_23763 & tmp_ivl_23758;
  tmp_ivl_23765 <= new_AGEMA_signal_3732 & n3828;
  LPM_q_ivl_23768 <= tmp_ivl_23770 & tmp_ivl_23765;
  new_AGEMA_signal_4056 <= tmp_ivl_23772(1);
  n3830 <= tmp_ivl_23772(0);
  tmp_ivl_23772 <= LPM_d0_ivl_23776(0 + 1 downto 0);
  tmp_ivl_23777 <= new_AGEMA_signal_4056 & n3830;
  LPM_q_ivl_23780 <= tmp_ivl_23782 & tmp_ivl_23777;
  tmp_ivl_23784 <= new_AGEMA_signal_3755 & n3829;
  LPM_q_ivl_23787 <= tmp_ivl_23789 & tmp_ivl_23784;
  tmp_ivl_23791 <= tmp_ivl_23795(1);
  tmp_ivl_23793 <= tmp_ivl_23795(0);
  tmp_ivl_23795 <= LPM_d0_ivl_23799(0 + 1 downto 0);
  tmp_ivl_23800 <= new_AGEMA_signal_3642 & n3832;
  LPM_q_ivl_23803 <= tmp_ivl_23805 & tmp_ivl_23800;
  tmp_ivl_23807 <= new_AGEMA_signal_3690 & n3831;
  LPM_q_ivl_23810 <= tmp_ivl_23812 & tmp_ivl_23807;
  new_AGEMA_signal_4057 <= tmp_ivl_23814(1);
  n3834 <= tmp_ivl_23814(0);
  tmp_ivl_23814 <= LPM_d0_ivl_23818(0 + 1 downto 0);
  tmp_ivl_23820 <= state_in_s1(267);
  tmp_ivl_23822 <= state_in_s0(267);
  tmp_ivl_23823 <= tmp_ivl_23820 & tmp_ivl_23822;
  LPM_q_ivl_23826 <= tmp_ivl_23828 & tmp_ivl_23823;
  tmp_ivl_23830 <= new_AGEMA_signal_3449 & n3833;
  LPM_q_ivl_23833 <= tmp_ivl_23835 & tmp_ivl_23830;
  new_AGEMA_signal_3756 <= tmp_ivl_23837(1);
  n3840 <= tmp_ivl_23837(0);
  tmp_ivl_23837 <= LPM_d0_ivl_23841(0 + 1 downto 0);
  tmp_ivl_23842 <= new_AGEMA_signal_4057 & n3834;
  LPM_q_ivl_23845 <= tmp_ivl_23847 & tmp_ivl_23842;
  tmp_ivl_23849 <= new_AGEMA_signal_3756 & n3840;
  LPM_q_ivl_23852 <= tmp_ivl_23854 & tmp_ivl_23849;
  tmp_ivl_23856 <= tmp_ivl_23860(1);
  tmp_ivl_23858 <= tmp_ivl_23860(0);
  tmp_ivl_23860 <= LPM_d0_ivl_23864(0 + 1 downto 0);
  tmp_ivl_23865 <= new_AGEMA_signal_3595 & n3836;
  LPM_q_ivl_23868 <= tmp_ivl_23870 & tmp_ivl_23865;
  tmp_ivl_23872 <= new_AGEMA_signal_3620 & n3835;
  LPM_q_ivl_23875 <= tmp_ivl_23877 & tmp_ivl_23872;
  new_AGEMA_signal_4058 <= tmp_ivl_23879(1);
  n3837 <= tmp_ivl_23879(0);
  tmp_ivl_23879 <= LPM_d0_ivl_23883(0 + 1 downto 0);
  tmp_ivl_23884 <= new_AGEMA_signal_4058 & n3837;
  LPM_q_ivl_23887 <= tmp_ivl_23889 & tmp_ivl_23884;
  tmp_ivl_23891 <= new_AGEMA_signal_3756 & n3840;
  LPM_q_ivl_23894 <= tmp_ivl_23896 & tmp_ivl_23891;
  tmp_ivl_23898 <= tmp_ivl_23902(1);
  tmp_ivl_23900 <= tmp_ivl_23902(0);
  tmp_ivl_23902 <= LPM_d0_ivl_23906(0 + 1 downto 0);
  tmp_ivl_23907 <= new_AGEMA_signal_3594 & n3839;
  LPM_q_ivl_23910 <= tmp_ivl_23912 & tmp_ivl_23907;
  tmp_ivl_23914 <= new_AGEMA_signal_3752 & n3838;
  LPM_q_ivl_23917 <= tmp_ivl_23919 & tmp_ivl_23914;
  new_AGEMA_signal_4059 <= tmp_ivl_23921(1);
  n3841 <= tmp_ivl_23921(0);
  tmp_ivl_23921 <= LPM_d0_ivl_23925(0 + 1 downto 0);
  tmp_ivl_23926 <= new_AGEMA_signal_4059 & n3841;
  LPM_q_ivl_23929 <= tmp_ivl_23931 & tmp_ivl_23926;
  tmp_ivl_23933 <= new_AGEMA_signal_3756 & n3840;
  LPM_q_ivl_23936 <= tmp_ivl_23938 & tmp_ivl_23933;
  tmp_ivl_23940 <= tmp_ivl_23944(1);
  tmp_ivl_23942 <= tmp_ivl_23944(0);
  tmp_ivl_23944 <= LPM_d0_ivl_23948(0 + 1 downto 0);
  tmp_ivl_23949 <= new_AGEMA_signal_3663 & n3843;
  LPM_q_ivl_23952 <= tmp_ivl_23954 & tmp_ivl_23949;
  tmp_ivl_23956 <= new_AGEMA_signal_4319 & n3842;
  LPM_q_ivl_23959 <= tmp_ivl_23961 & tmp_ivl_23956;
  new_AGEMA_signal_4511 <= tmp_ivl_23963(1);
  n3845 <= tmp_ivl_23963(0);
  tmp_ivl_23963 <= LPM_d0_ivl_23967(0 + 1 downto 0);
  tmp_ivl_23969 <= z0(46);
  tmp_ivl_23970 <= new_AGEMA_signal_3213 & tmp_ivl_23969;
  LPM_q_ivl_23973 <= tmp_ivl_23975 & tmp_ivl_23970;
  tmp_ivl_23978 <= state_in_s1(22);
  tmp_ivl_23980 <= state_in_s0(22);
  tmp_ivl_23981 <= tmp_ivl_23978 & tmp_ivl_23980;
  LPM_q_ivl_23984 <= tmp_ivl_23986 & tmp_ivl_23981;
  new_AGEMA_signal_3450 <= tmp_ivl_23988(1);
  n3849 <= tmp_ivl_23988(0);
  tmp_ivl_23988 <= LPM_d0_ivl_23992(0 + 1 downto 0);
  tmp_ivl_23993 <= new_AGEMA_signal_3450 & n3849;
  LPM_q_ivl_23996 <= tmp_ivl_23998 & tmp_ivl_23993;
  tmp_ivl_24000 <= new_AGEMA_signal_3313 & n3844;
  LPM_q_ivl_24003 <= tmp_ivl_24005 & tmp_ivl_24000;
  new_AGEMA_signal_3757 <= tmp_ivl_24007(1);
  n3862 <= tmp_ivl_24007(0);
  tmp_ivl_24007 <= LPM_d0_ivl_24011(0 + 1 downto 0);
  tmp_ivl_24012 <= new_AGEMA_signal_4511 & n3845;
  LPM_q_ivl_24015 <= tmp_ivl_24017 & tmp_ivl_24012;
  tmp_ivl_24019 <= new_AGEMA_signal_3757 & n3862;
  LPM_q_ivl_24022 <= tmp_ivl_24024 & tmp_ivl_24019;
  tmp_ivl_24026 <= tmp_ivl_24030(1);
  tmp_ivl_24028 <= tmp_ivl_24030(0);
  tmp_ivl_24030 <= LPM_d0_ivl_24034(0 + 1 downto 0);
  tmp_ivl_24035 <= new_AGEMA_signal_3662 & n3846;
  LPM_q_ivl_24038 <= tmp_ivl_24040 & tmp_ivl_24035;
  tmp_ivl_24042 <= new_AGEMA_signal_3671 & n3856;
  LPM_q_ivl_24045 <= tmp_ivl_24047 & tmp_ivl_24042;
  new_AGEMA_signal_4060 <= tmp_ivl_24049(1);
  n3847 <= tmp_ivl_24049(0);
  tmp_ivl_24049 <= LPM_d0_ivl_24053(0 + 1 downto 0);
  tmp_ivl_24054 <= new_AGEMA_signal_4060 & n3847;
  LPM_q_ivl_24057 <= tmp_ivl_24059 & tmp_ivl_24054;
  tmp_ivl_24061 <= new_AGEMA_signal_3757 & n3862;
  LPM_q_ivl_24064 <= tmp_ivl_24066 & tmp_ivl_24061;
  tmp_ivl_24068 <= tmp_ivl_24072(1);
  tmp_ivl_24070 <= tmp_ivl_24072(0);
  tmp_ivl_24072 <= LPM_d0_ivl_24076(0 + 1 downto 0);
  tmp_ivl_24077 <= new_AGEMA_signal_3955 & n3883;
  LPM_q_ivl_24080 <= tmp_ivl_24082 & tmp_ivl_24077;
  tmp_ivl_24084 <= new_AGEMA_signal_3997 & n3848;
  LPM_q_ivl_24087 <= tmp_ivl_24089 & tmp_ivl_24084;
  new_AGEMA_signal_4364 <= tmp_ivl_24091(1);
  n3852 <= tmp_ivl_24091(0);
  tmp_ivl_24091 <= LPM_d0_ivl_24095(0 + 1 downto 0);
  tmp_ivl_24097 <= z1(46);
  tmp_ivl_24098 <= new_AGEMA_signal_3027 & tmp_ivl_24097;
  LPM_q_ivl_24101 <= tmp_ivl_24103 & tmp_ivl_24098;
  tmp_ivl_24106 <= state_in_s1(278);
  tmp_ivl_24108 <= state_in_s0(278);
  tmp_ivl_24109 <= tmp_ivl_24106 & tmp_ivl_24108;
  LPM_q_ivl_24112 <= tmp_ivl_24114 & tmp_ivl_24109;
  new_AGEMA_signal_3451 <= tmp_ivl_24116(1);
  n3851 <= tmp_ivl_24116(0);
  tmp_ivl_24116 <= LPM_d0_ivl_24120(0 + 1 downto 0);
  tmp_ivl_24122 <= state_in_s1(86);
  tmp_ivl_24124 <= state_in_s0(86);
  tmp_ivl_24125 <= tmp_ivl_24122 & tmp_ivl_24124;
  LPM_q_ivl_24128 <= tmp_ivl_24130 & tmp_ivl_24125;
  tmp_ivl_24132 <= new_AGEMA_signal_3450 & n3849;
  LPM_q_ivl_24135 <= tmp_ivl_24137 & tmp_ivl_24132;
  new_AGEMA_signal_3758 <= tmp_ivl_24139(1);
  n3850 <= tmp_ivl_24139(0);
  tmp_ivl_24139 <= LPM_d0_ivl_24143(0 + 1 downto 0);
  tmp_ivl_24144 <= new_AGEMA_signal_3451 & n3851;
  LPM_q_ivl_24147 <= tmp_ivl_24149 & tmp_ivl_24144;
  tmp_ivl_24151 <= new_AGEMA_signal_3758 & n3850;
  LPM_q_ivl_24154 <= tmp_ivl_24156 & tmp_ivl_24151;
  new_AGEMA_signal_4061 <= tmp_ivl_24158(1);
  n3907 <= tmp_ivl_24158(0);
  tmp_ivl_24158 <= LPM_d0_ivl_24162(0 + 1 downto 0);
  tmp_ivl_24163 <= new_AGEMA_signal_4364 & n3852;
  LPM_q_ivl_24166 <= tmp_ivl_24168 & tmp_ivl_24163;
  tmp_ivl_24170 <= new_AGEMA_signal_4061 & n3907;
  LPM_q_ivl_24173 <= tmp_ivl_24175 & tmp_ivl_24170;
  tmp_ivl_24177 <= tmp_ivl_24181(1);
  tmp_ivl_24179 <= tmp_ivl_24181(0);
  tmp_ivl_24181 <= LPM_d0_ivl_24185(0 + 1 downto 0);
  tmp_ivl_24186 <= new_AGEMA_signal_3919 & n3853;
  LPM_q_ivl_24189 <= tmp_ivl_24191 & tmp_ivl_24186;
  tmp_ivl_24193 <= new_AGEMA_signal_4013 & n3904;
  LPM_q_ivl_24196 <= tmp_ivl_24198 & tmp_ivl_24193;
  new_AGEMA_signal_4365 <= tmp_ivl_24200(1);
  n3854 <= tmp_ivl_24200(0);
  tmp_ivl_24200 <= LPM_d0_ivl_24204(0 + 1 downto 0);
  tmp_ivl_24205 <= new_AGEMA_signal_4365 & n3854;
  LPM_q_ivl_24208 <= tmp_ivl_24210 & tmp_ivl_24205;
  tmp_ivl_24212 <= new_AGEMA_signal_4061 & n3907;
  LPM_q_ivl_24215 <= tmp_ivl_24217 & tmp_ivl_24212;
  tmp_ivl_24219 <= tmp_ivl_24223(1);
  tmp_ivl_24221 <= tmp_ivl_24223(0);
  tmp_ivl_24223 <= LPM_d0_ivl_24227(0 + 1 downto 0);
  tmp_ivl_24228 <= new_AGEMA_signal_3671 & n3856;
  LPM_q_ivl_24231 <= tmp_ivl_24233 & tmp_ivl_24228;
  tmp_ivl_24235 <= new_AGEMA_signal_3721 & n3855;
  LPM_q_ivl_24238 <= tmp_ivl_24240 & tmp_ivl_24235;
  new_AGEMA_signal_4062 <= tmp_ivl_24242(1);
  n3858 <= tmp_ivl_24242(0);
  tmp_ivl_24242 <= LPM_d0_ivl_24246(0 + 1 downto 0);
  tmp_ivl_24248 <= state_in_s1(234);
  tmp_ivl_24250 <= state_in_s0(234);
  tmp_ivl_24251 <= tmp_ivl_24248 & tmp_ivl_24250;
  LPM_q_ivl_24254 <= tmp_ivl_24256 & tmp_ivl_24251;
  tmp_ivl_24259 <= z4(18);
  tmp_ivl_24260 <= new_AGEMA_signal_3120 & tmp_ivl_24259;
  LPM_q_ivl_24263 <= tmp_ivl_24265 & tmp_ivl_24260;
  new_AGEMA_signal_3452 <= tmp_ivl_24267(1);
  n3868 <= tmp_ivl_24267(0);
  tmp_ivl_24267 <= LPM_d0_ivl_24271(0 + 1 downto 0);
  tmp_ivl_24272 <= new_AGEMA_signal_3353 & n3857;
  LPM_q_ivl_24275 <= tmp_ivl_24277 & tmp_ivl_24272;
  tmp_ivl_24279 <= new_AGEMA_signal_3452 & n3868;
  LPM_q_ivl_24282 <= tmp_ivl_24284 & tmp_ivl_24279;
  new_AGEMA_signal_3759 <= tmp_ivl_24286(1);
  n3864 <= tmp_ivl_24286(0);
  tmp_ivl_24286 <= LPM_d0_ivl_24290(0 + 1 downto 0);
  tmp_ivl_24291 <= new_AGEMA_signal_4062 & n3858;
  LPM_q_ivl_24294 <= tmp_ivl_24296 & tmp_ivl_24291;
  tmp_ivl_24298 <= new_AGEMA_signal_3759 & n3864;
  LPM_q_ivl_24301 <= tmp_ivl_24303 & tmp_ivl_24298;
  tmp_ivl_24305 <= tmp_ivl_24309(1);
  tmp_ivl_24307 <= tmp_ivl_24309(0);
  tmp_ivl_24309 <= LPM_d0_ivl_24313(0 + 1 downto 0);
  tmp_ivl_24314 <= new_AGEMA_signal_3689 & n3860;
  LPM_q_ivl_24317 <= tmp_ivl_24319 & tmp_ivl_24314;
  tmp_ivl_24321 <= new_AGEMA_signal_3720 & n3859;
  LPM_q_ivl_24324 <= tmp_ivl_24326 & tmp_ivl_24321;
  new_AGEMA_signal_4063 <= tmp_ivl_24328(1);
  n3861 <= tmp_ivl_24328(0);
  tmp_ivl_24328 <= LPM_d0_ivl_24332(0 + 1 downto 0);
  tmp_ivl_24333 <= new_AGEMA_signal_4063 & n3861;
  LPM_q_ivl_24336 <= tmp_ivl_24338 & tmp_ivl_24333;
  tmp_ivl_24340 <= new_AGEMA_signal_3759 & n3864;
  LPM_q_ivl_24343 <= tmp_ivl_24345 & tmp_ivl_24340;
  tmp_ivl_24347 <= tmp_ivl_24351(1);
  tmp_ivl_24349 <= tmp_ivl_24351(0);
  tmp_ivl_24351 <= LPM_d0_ivl_24355(0 + 1 downto 0);
  tmp_ivl_24356 <= new_AGEMA_signal_3688 & n3863;
  LPM_q_ivl_24359 <= tmp_ivl_24361 & tmp_ivl_24356;
  tmp_ivl_24363 <= new_AGEMA_signal_3757 & n3862;
  LPM_q_ivl_24366 <= tmp_ivl_24368 & tmp_ivl_24363;
  new_AGEMA_signal_4064 <= tmp_ivl_24370(1);
  n3865 <= tmp_ivl_24370(0);
  tmp_ivl_24370 <= LPM_d0_ivl_24374(0 + 1 downto 0);
  tmp_ivl_24375 <= new_AGEMA_signal_4064 & n3865;
  LPM_q_ivl_24378 <= tmp_ivl_24380 & tmp_ivl_24375;
  tmp_ivl_24382 <= new_AGEMA_signal_3759 & n3864;
  LPM_q_ivl_24385 <= tmp_ivl_24387 & tmp_ivl_24382;
  tmp_ivl_24389 <= tmp_ivl_24393(1);
  tmp_ivl_24391 <= tmp_ivl_24393(0);
  tmp_ivl_24393 <= LPM_d0_ivl_24397(0 + 1 downto 0);
  tmp_ivl_24398 <= new_AGEMA_signal_3614 & n3867;
  LPM_q_ivl_24401 <= tmp_ivl_24403 & tmp_ivl_24398;
  tmp_ivl_24405 <= new_AGEMA_signal_3647 & n3866;
  LPM_q_ivl_24408 <= tmp_ivl_24410 & tmp_ivl_24405;
  new_AGEMA_signal_4065 <= tmp_ivl_24412(1);
  n3869 <= tmp_ivl_24412(0);
  tmp_ivl_24412 <= LPM_d0_ivl_24416(0 + 1 downto 0);
  tmp_ivl_24418 <= state_in_s1(298);
  tmp_ivl_24420 <= state_in_s0(298);
  tmp_ivl_24421 <= tmp_ivl_24418 & tmp_ivl_24420;
  LPM_q_ivl_24424 <= tmp_ivl_24426 & tmp_ivl_24421;
  tmp_ivl_24428 <= new_AGEMA_signal_3452 & n3868;
  LPM_q_ivl_24431 <= tmp_ivl_24433 & tmp_ivl_24428;
  new_AGEMA_signal_3760 <= tmp_ivl_24435(1);
  n3928 <= tmp_ivl_24435(0);
  tmp_ivl_24435 <= LPM_d0_ivl_24439(0 + 1 downto 0);
  tmp_ivl_24440 <= new_AGEMA_signal_4065 & n3869;
  LPM_q_ivl_24443 <= tmp_ivl_24445 & tmp_ivl_24440;
  tmp_ivl_24447 <= new_AGEMA_signal_3760 & n3928;
  LPM_q_ivl_24450 <= tmp_ivl_24452 & tmp_ivl_24447;
  tmp_ivl_24454 <= tmp_ivl_24458(1);
  tmp_ivl_24456 <= tmp_ivl_24458(0);
  tmp_ivl_24458 <= LPM_d0_ivl_24462(0 + 1 downto 0);
  tmp_ivl_24463 <= new_AGEMA_signal_3646 & n3870;
  LPM_q_ivl_24466 <= tmp_ivl_24468 & tmp_ivl_24463;
  tmp_ivl_24470 <= new_AGEMA_signal_3648 & n3922;
  LPM_q_ivl_24473 <= tmp_ivl_24475 & tmp_ivl_24470;
  new_AGEMA_signal_4066 <= tmp_ivl_24477(1);
  n3871 <= tmp_ivl_24477(0);
  tmp_ivl_24477 <= LPM_d0_ivl_24481(0 + 1 downto 0);
  tmp_ivl_24482 <= new_AGEMA_signal_4066 & n3871;
  LPM_q_ivl_24485 <= tmp_ivl_24487 & tmp_ivl_24482;
  tmp_ivl_24489 <= new_AGEMA_signal_3760 & n3928;
  LPM_q_ivl_24492 <= tmp_ivl_24494 & tmp_ivl_24489;
  tmp_ivl_24496 <= tmp_ivl_24500(1);
  tmp_ivl_24498 <= tmp_ivl_24500(0);
  tmp_ivl_24500 <= LPM_d0_ivl_24504(0 + 1 downto 0);
  tmp_ivl_24505 <= new_AGEMA_signal_3714 & n3872;
  LPM_q_ivl_24508 <= tmp_ivl_24510 & tmp_ivl_24505;
  tmp_ivl_24512 <= new_AGEMA_signal_3738 & n3917;
  LPM_q_ivl_24515 <= tmp_ivl_24517 & tmp_ivl_24512;
  new_AGEMA_signal_4067 <= tmp_ivl_24519(1);
  n3874 <= tmp_ivl_24519(0);
  tmp_ivl_24519 <= LPM_d0_ivl_24523(0 + 1 downto 0);
  tmp_ivl_24525 <= z0(7);
  tmp_ivl_24526 <= new_AGEMA_signal_4579 & tmp_ivl_24525;
  LPM_q_ivl_24529 <= tmp_ivl_24531 & tmp_ivl_24526;
  tmp_ivl_24534 <= state_in_s1(63);
  tmp_ivl_24536 <= state_in_s0(63);
  tmp_ivl_24537 <= tmp_ivl_24534 & tmp_ivl_24536;
  LPM_q_ivl_24540 <= tmp_ivl_24542 & tmp_ivl_24537;
  new_AGEMA_signal_4596 <= tmp_ivl_24544(1);
  n3879 <= tmp_ivl_24544(0);
  tmp_ivl_24544 <= LPM_d0_ivl_24548(0 + 1 downto 0);
  tmp_ivl_24549 <= new_AGEMA_signal_4596 & n3879;
  LPM_q_ivl_24552 <= tmp_ivl_24554 & tmp_ivl_24549;
  tmp_ivl_24556 <= new_AGEMA_signal_3376 & n3873;
  LPM_q_ivl_24559 <= tmp_ivl_24561 & tmp_ivl_24556;
  new_AGEMA_signal_4621 <= tmp_ivl_24563(1);
  n3910 <= tmp_ivl_24563(0);
  tmp_ivl_24563 <= LPM_d0_ivl_24567(0 + 1 downto 0);
  tmp_ivl_24568 <= new_AGEMA_signal_4067 & n3874;
  LPM_q_ivl_24571 <= tmp_ivl_24573 & tmp_ivl_24568;
  tmp_ivl_24575 <= new_AGEMA_signal_4621 & n3910;
  LPM_q_ivl_24578 <= tmp_ivl_24580 & tmp_ivl_24575;
  tmp_ivl_24582 <= tmp_ivl_24586(1);
  tmp_ivl_24584 <= tmp_ivl_24586(0);
  tmp_ivl_24586 <= LPM_d0_ivl_24590(0 + 1 downto 0);
  tmp_ivl_24591 <= new_AGEMA_signal_3719 & n3876;
  LPM_q_ivl_24594 <= tmp_ivl_24596 & tmp_ivl_24591;
  tmp_ivl_24598 <= new_AGEMA_signal_3750 & n3875;
  LPM_q_ivl_24601 <= tmp_ivl_24603 & tmp_ivl_24598;
  new_AGEMA_signal_4068 <= tmp_ivl_24605(1);
  n3877 <= tmp_ivl_24605(0);
  tmp_ivl_24605 <= LPM_d0_ivl_24609(0 + 1 downto 0);
  tmp_ivl_24610 <= new_AGEMA_signal_4068 & n3877;
  LPM_q_ivl_24613 <= tmp_ivl_24615 & tmp_ivl_24610;
  tmp_ivl_24617 <= new_AGEMA_signal_4621 & n3910;
  LPM_q_ivl_24620 <= tmp_ivl_24622 & tmp_ivl_24617;
  tmp_ivl_24624 <= tmp_ivl_24628(1);
  tmp_ivl_24626 <= tmp_ivl_24628(0);
  tmp_ivl_24628 <= LPM_d0_ivl_24632(0 + 1 downto 0);
  tmp_ivl_24633 <= new_AGEMA_signal_3949 & n3878;
  LPM_q_ivl_24636 <= tmp_ivl_24638 & tmp_ivl_24633;
  tmp_ivl_24640 <= new_AGEMA_signal_3979 & n3897;
  LPM_q_ivl_24643 <= tmp_ivl_24645 & tmp_ivl_24640;
  new_AGEMA_signal_4371 <= tmp_ivl_24647(1);
  n3882 <= tmp_ivl_24647(0);
  tmp_ivl_24647 <= LPM_d0_ivl_24651(0 + 1 downto 0);
  tmp_ivl_24653 <= z1(7);
  tmp_ivl_24654 <= new_AGEMA_signal_4578 & tmp_ivl_24653;
  LPM_q_ivl_24657 <= tmp_ivl_24659 & tmp_ivl_24654;
  tmp_ivl_24662 <= state_in_s1(319);
  tmp_ivl_24664 <= state_in_s0(319);
  tmp_ivl_24665 <= tmp_ivl_24662 & tmp_ivl_24664;
  LPM_q_ivl_24668 <= tmp_ivl_24670 & tmp_ivl_24665;
  new_AGEMA_signal_4597 <= tmp_ivl_24672(1);
  n3881 <= tmp_ivl_24672(0);
  tmp_ivl_24672 <= LPM_d0_ivl_24676(0 + 1 downto 0);
  tmp_ivl_24678 <= state_in_s1(127);
  tmp_ivl_24680 <= state_in_s0(127);
  tmp_ivl_24681 <= tmp_ivl_24678 & tmp_ivl_24680;
  LPM_q_ivl_24684 <= tmp_ivl_24686 & tmp_ivl_24681;
  tmp_ivl_24688 <= new_AGEMA_signal_4596 & n3879;
  LPM_q_ivl_24691 <= tmp_ivl_24693 & tmp_ivl_24688;
  new_AGEMA_signal_4622 <= tmp_ivl_24695(1);
  n3880 <= tmp_ivl_24695(0);
  tmp_ivl_24695 <= LPM_d0_ivl_24699(0 + 1 downto 0);
  tmp_ivl_24700 <= new_AGEMA_signal_4597 & n3881;
  LPM_q_ivl_24703 <= tmp_ivl_24705 & tmp_ivl_24700;
  tmp_ivl_24707 <= new_AGEMA_signal_4622 & n3880;
  LPM_q_ivl_24710 <= tmp_ivl_24712 & tmp_ivl_24707;
  new_AGEMA_signal_4642 <= tmp_ivl_24714(1);
  n3906 <= tmp_ivl_24714(0);
  tmp_ivl_24714 <= LPM_d0_ivl_24718(0 + 1 downto 0);
  tmp_ivl_24719 <= new_AGEMA_signal_4371 & n3882;
  LPM_q_ivl_24722 <= tmp_ivl_24724 & tmp_ivl_24719;
  tmp_ivl_24726 <= new_AGEMA_signal_4642 & n3906;
  LPM_q_ivl_24729 <= tmp_ivl_24731 & tmp_ivl_24726;
  tmp_ivl_24733 <= tmp_ivl_24737(1);
  tmp_ivl_24735 <= tmp_ivl_24737(0);
  tmp_ivl_24737 <= LPM_d0_ivl_24741(0 + 1 downto 0);
  tmp_ivl_24742 <= new_AGEMA_signal_3948 & n3884;
  LPM_q_ivl_24745 <= tmp_ivl_24747 & tmp_ivl_24742;
  tmp_ivl_24749 <= new_AGEMA_signal_3955 & n3883;
  LPM_q_ivl_24752 <= tmp_ivl_24754 & tmp_ivl_24749;
  new_AGEMA_signal_4372 <= tmp_ivl_24756(1);
  n3885 <= tmp_ivl_24756(0);
  tmp_ivl_24756 <= LPM_d0_ivl_24760(0 + 1 downto 0);
  tmp_ivl_24761 <= new_AGEMA_signal_4372 & n3885;
  LPM_q_ivl_24764 <= tmp_ivl_24766 & tmp_ivl_24761;
  tmp_ivl_24768 <= new_AGEMA_signal_4642 & n3906;
  LPM_q_ivl_24771 <= tmp_ivl_24773 & tmp_ivl_24768;
  tmp_ivl_24775 <= tmp_ivl_24779(1);
  tmp_ivl_24777 <= tmp_ivl_24779(0);
  tmp_ivl_24779 <= LPM_d0_ivl_24783(0 + 1 downto 0);
  tmp_ivl_24784 <= new_AGEMA_signal_3666 & n3887;
  LPM_q_ivl_24787 <= tmp_ivl_24789 & tmp_ivl_24784;
  tmp_ivl_24791 <= new_AGEMA_signal_3740 & n3886;
  LPM_q_ivl_24794 <= tmp_ivl_24796 & tmp_ivl_24791;
  new_AGEMA_signal_4069 <= tmp_ivl_24798(1);
  n3889 <= tmp_ivl_24798(0);
  tmp_ivl_24798 <= LPM_d0_ivl_24802(0 + 1 downto 0);
  tmp_ivl_24804 <= z0(4);
  tmp_ivl_24805 <= new_AGEMA_signal_3583 & tmp_ivl_24804;
  LPM_q_ivl_24808 <= tmp_ivl_24810 & tmp_ivl_24805;
  tmp_ivl_24813 <= state_in_s1(60);
  tmp_ivl_24815 <= state_in_s0(60);
  tmp_ivl_24816 <= tmp_ivl_24813 & tmp_ivl_24815;
  LPM_q_ivl_24819 <= tmp_ivl_24821 & tmp_ivl_24816;
  new_AGEMA_signal_3761 <= tmp_ivl_24823(1);
  n3899 <= tmp_ivl_24823(0);
  tmp_ivl_24823 <= LPM_d0_ivl_24827(0 + 1 downto 0);
  tmp_ivl_24828 <= new_AGEMA_signal_3761 & n3899;
  LPM_q_ivl_24831 <= tmp_ivl_24833 & tmp_ivl_24828;
  tmp_ivl_24835 <= new_AGEMA_signal_3309 & n3888;
  LPM_q_ivl_24838 <= tmp_ivl_24840 & tmp_ivl_24835;
  new_AGEMA_signal_4070 <= tmp_ivl_24842(1);
  n3895 <= tmp_ivl_24842(0);
  tmp_ivl_24842 <= LPM_d0_ivl_24846(0 + 1 downto 0);
  tmp_ivl_24847 <= new_AGEMA_signal_4069 & n3889;
  LPM_q_ivl_24850 <= tmp_ivl_24852 & tmp_ivl_24847;
  tmp_ivl_24854 <= new_AGEMA_signal_4070 & n3895;
  LPM_q_ivl_24857 <= tmp_ivl_24859 & tmp_ivl_24854;
  tmp_ivl_24861 <= tmp_ivl_24865(1);
  tmp_ivl_24863 <= tmp_ivl_24865(0);
  tmp_ivl_24865 <= LPM_d0_ivl_24869(0 + 1 downto 0);
  tmp_ivl_24870 <= new_AGEMA_signal_3710 & n3891;
  LPM_q_ivl_24873 <= tmp_ivl_24875 & tmp_ivl_24870;
  tmp_ivl_24877 <= new_AGEMA_signal_3725 & n3890;
  LPM_q_ivl_24880 <= tmp_ivl_24882 & tmp_ivl_24877;
  new_AGEMA_signal_4071 <= tmp_ivl_24884(1);
  n3892 <= tmp_ivl_24884(0);
  tmp_ivl_24884 <= LPM_d0_ivl_24888(0 + 1 downto 0);
  tmp_ivl_24889 <= new_AGEMA_signal_4071 & n3892;
  LPM_q_ivl_24892 <= tmp_ivl_24894 & tmp_ivl_24889;
  tmp_ivl_24896 <= new_AGEMA_signal_4070 & n3895;
  LPM_q_ivl_24899 <= tmp_ivl_24901 & tmp_ivl_24896;
  tmp_ivl_24903 <= tmp_ivl_24907(1);
  tmp_ivl_24905 <= tmp_ivl_24907(0);
  tmp_ivl_24907 <= LPM_d0_ivl_24911(0 + 1 downto 0);
  tmp_ivl_24912 <= new_AGEMA_signal_3724 & n3894;
  LPM_q_ivl_24915 <= tmp_ivl_24917 & tmp_ivl_24912;
  tmp_ivl_24919 <= new_AGEMA_signal_3728 & n3893;
  LPM_q_ivl_24922 <= tmp_ivl_24924 & tmp_ivl_24919;
  new_AGEMA_signal_4072 <= tmp_ivl_24926(1);
  n3896 <= tmp_ivl_24926(0);
  tmp_ivl_24926 <= LPM_d0_ivl_24930(0 + 1 downto 0);
  tmp_ivl_24931 <= new_AGEMA_signal_4072 & n3896;
  LPM_q_ivl_24934 <= tmp_ivl_24936 & tmp_ivl_24931;
  tmp_ivl_24938 <= new_AGEMA_signal_4070 & n3895;
  LPM_q_ivl_24941 <= tmp_ivl_24943 & tmp_ivl_24938;
  tmp_ivl_24945 <= tmp_ivl_24949(1);
  tmp_ivl_24947 <= tmp_ivl_24949(0);
  tmp_ivl_24949 <= LPM_d0_ivl_24953(0 + 1 downto 0);
  tmp_ivl_24954 <= new_AGEMA_signal_3942 & n3898;
  LPM_q_ivl_24957 <= tmp_ivl_24959 & tmp_ivl_24954;
  tmp_ivl_24961 <= new_AGEMA_signal_3979 & n3897;
  LPM_q_ivl_24964 <= tmp_ivl_24966 & tmp_ivl_24961;
  new_AGEMA_signal_4376 <= tmp_ivl_24968(1);
  n3902 <= tmp_ivl_24968(0);
  tmp_ivl_24968 <= LPM_d0_ivl_24972(0 + 1 downto 0);
  tmp_ivl_24974 <= z1(4);
  tmp_ivl_24975 <= new_AGEMA_signal_3518 & tmp_ivl_24974;
  LPM_q_ivl_24978 <= tmp_ivl_24980 & tmp_ivl_24975;
  tmp_ivl_24983 <= state_in_s1(316);
  tmp_ivl_24985 <= state_in_s0(316);
  tmp_ivl_24986 <= tmp_ivl_24983 & tmp_ivl_24985;
  LPM_q_ivl_24989 <= tmp_ivl_24991 & tmp_ivl_24986;
  new_AGEMA_signal_3762 <= tmp_ivl_24993(1);
  n3901 <= tmp_ivl_24993(0);
  tmp_ivl_24993 <= LPM_d0_ivl_24997(0 + 1 downto 0);
  tmp_ivl_24999 <= state_in_s1(124);
  tmp_ivl_25001 <= state_in_s0(124);
  tmp_ivl_25002 <= tmp_ivl_24999 & tmp_ivl_25001;
  LPM_q_ivl_25005 <= tmp_ivl_25007 & tmp_ivl_25002;
  tmp_ivl_25009 <= new_AGEMA_signal_3761 & n3899;
  LPM_q_ivl_25012 <= tmp_ivl_25014 & tmp_ivl_25009;
  new_AGEMA_signal_4073 <= tmp_ivl_25016(1);
  n3900 <= tmp_ivl_25016(0);
  tmp_ivl_25016 <= LPM_d0_ivl_25020(0 + 1 downto 0);
  tmp_ivl_25021 <= new_AGEMA_signal_3762 & n3901;
  LPM_q_ivl_25024 <= tmp_ivl_25026 & tmp_ivl_25021;
  tmp_ivl_25028 <= new_AGEMA_signal_4073 & n3900;
  LPM_q_ivl_25031 <= tmp_ivl_25033 & tmp_ivl_25028;
  new_AGEMA_signal_4377 <= tmp_ivl_25035(1);
  n3908 <= tmp_ivl_25035(0);
  tmp_ivl_25035 <= LPM_d0_ivl_25039(0 + 1 downto 0);
  tmp_ivl_25040 <= new_AGEMA_signal_4376 & n3902;
  LPM_q_ivl_25043 <= tmp_ivl_25045 & tmp_ivl_25040;
  tmp_ivl_25047 <= new_AGEMA_signal_4377 & n3908;
  LPM_q_ivl_25050 <= tmp_ivl_25052 & tmp_ivl_25047;
  tmp_ivl_25054 <= tmp_ivl_25058(1);
  tmp_ivl_25056 <= tmp_ivl_25058(0);
  tmp_ivl_25058 <= LPM_d0_ivl_25062(0 + 1 downto 0);
  tmp_ivl_25063 <= new_AGEMA_signal_4013 & n3904;
  LPM_q_ivl_25066 <= tmp_ivl_25068 & tmp_ivl_25063;
  tmp_ivl_25070 <= new_AGEMA_signal_4496 & n3903;
  LPM_q_ivl_25073 <= tmp_ivl_25075 & tmp_ivl_25070;
  new_AGEMA_signal_4598 <= tmp_ivl_25077(1);
  n3905 <= tmp_ivl_25077(0);
  tmp_ivl_25077 <= LPM_d0_ivl_25081(0 + 1 downto 0);
  tmp_ivl_25082 <= new_AGEMA_signal_4598 & n3905;
  LPM_q_ivl_25085 <= tmp_ivl_25087 & tmp_ivl_25082;
  tmp_ivl_25089 <= new_AGEMA_signal_4377 & n3908;
  LPM_q_ivl_25092 <= tmp_ivl_25094 & tmp_ivl_25089;
  tmp_ivl_25096 <= tmp_ivl_25100(1);
  tmp_ivl_25098 <= tmp_ivl_25100(0);
  tmp_ivl_25100 <= LPM_d0_ivl_25104(0 + 1 downto 0);
  tmp_ivl_25105 <= new_AGEMA_signal_4061 & n3907;
  LPM_q_ivl_25108 <= tmp_ivl_25110 & tmp_ivl_25105;
  tmp_ivl_25112 <= new_AGEMA_signal_4642 & n3906;
  LPM_q_ivl_25115 <= tmp_ivl_25117 & tmp_ivl_25112;
  new_AGEMA_signal_4651 <= tmp_ivl_25119(1);
  n3909 <= tmp_ivl_25119(0);
  tmp_ivl_25119 <= LPM_d0_ivl_25123(0 + 1 downto 0);
  tmp_ivl_25124 <= new_AGEMA_signal_4651 & n3909;
  LPM_q_ivl_25127 <= tmp_ivl_25129 & tmp_ivl_25124;
  tmp_ivl_25131 <= new_AGEMA_signal_4377 & n3908;
  LPM_q_ivl_25134 <= tmp_ivl_25136 & tmp_ivl_25131;
  tmp_ivl_25138 <= tmp_ivl_25142(1);
  tmp_ivl_25140 <= tmp_ivl_25142(0);
  tmp_ivl_25142 <= LPM_d0_ivl_25146(0 + 1 downto 0);
  tmp_ivl_25147 <= new_AGEMA_signal_3743 & n3911;
  LPM_q_ivl_25150 <= tmp_ivl_25152 & tmp_ivl_25147;
  tmp_ivl_25154 <= new_AGEMA_signal_4621 & n3910;
  LPM_q_ivl_25157 <= tmp_ivl_25159 & tmp_ivl_25154;
  new_AGEMA_signal_4643 <= tmp_ivl_25161(1);
  n3913 <= tmp_ivl_25161(0);
  tmp_ivl_25161 <= LPM_d0_ivl_25165(0 + 1 downto 0);
  tmp_ivl_25167 <= state_in_s1(204);
  tmp_ivl_25169 <= state_in_s0(204);
  tmp_ivl_25170 <= tmp_ivl_25167 & tmp_ivl_25169;
  LPM_q_ivl_25173 <= tmp_ivl_25175 & tmp_ivl_25170;
  tmp_ivl_25178 <= z4(52);
  tmp_ivl_25179 <= new_AGEMA_signal_3158 & tmp_ivl_25178;
  LPM_q_ivl_25182 <= tmp_ivl_25184 & tmp_ivl_25179;
  new_AGEMA_signal_3453 <= tmp_ivl_25186(1);
  n3923 <= tmp_ivl_25186(0);
  tmp_ivl_25186 <= LPM_d0_ivl_25190(0 + 1 downto 0);
  tmp_ivl_25191 <= new_AGEMA_signal_3400 & n3912;
  LPM_q_ivl_25194 <= tmp_ivl_25196 & tmp_ivl_25191;
  tmp_ivl_25198 <= new_AGEMA_signal_3453 & n3923;
  LPM_q_ivl_25201 <= tmp_ivl_25203 & tmp_ivl_25198;
  new_AGEMA_signal_3763 <= tmp_ivl_25205(1);
  n3919 <= tmp_ivl_25205(0);
  tmp_ivl_25205 <= LPM_d0_ivl_25209(0 + 1 downto 0);
  tmp_ivl_25210 <= new_AGEMA_signal_4643 & n3913;
  LPM_q_ivl_25213 <= tmp_ivl_25215 & tmp_ivl_25210;
  tmp_ivl_25217 <= new_AGEMA_signal_3763 & n3919;
  LPM_q_ivl_25220 <= tmp_ivl_25222 & tmp_ivl_25217;
  tmp_ivl_25224 <= tmp_ivl_25228(1);
  tmp_ivl_25226 <= tmp_ivl_25228(0);
  tmp_ivl_25228 <= LPM_d0_ivl_25232(0 + 1 downto 0);
  tmp_ivl_25233 <= new_AGEMA_signal_3731 & n3915;
  LPM_q_ivl_25236 <= tmp_ivl_25238 & tmp_ivl_25233;
  tmp_ivl_25240 <= new_AGEMA_signal_3742 & n3914;
  LPM_q_ivl_25243 <= tmp_ivl_25245 & tmp_ivl_25240;
  new_AGEMA_signal_4074 <= tmp_ivl_25247(1);
  n3916 <= tmp_ivl_25247(0);
  tmp_ivl_25247 <= LPM_d0_ivl_25251(0 + 1 downto 0);
  tmp_ivl_25252 <= new_AGEMA_signal_4074 & n3916;
  LPM_q_ivl_25255 <= tmp_ivl_25257 & tmp_ivl_25252;
  tmp_ivl_25259 <= new_AGEMA_signal_3763 & n3919;
  LPM_q_ivl_25262 <= tmp_ivl_25264 & tmp_ivl_25259;
  tmp_ivl_25266 <= tmp_ivl_25270(1);
  tmp_ivl_25268 <= tmp_ivl_25270(0);
  tmp_ivl_25270 <= LPM_d0_ivl_25274(0 + 1 downto 0);
  tmp_ivl_25275 <= new_AGEMA_signal_3691 & n3918;
  LPM_q_ivl_25278 <= tmp_ivl_25280 & tmp_ivl_25275;
  tmp_ivl_25282 <= new_AGEMA_signal_3738 & n3917;
  LPM_q_ivl_25285 <= tmp_ivl_25287 & tmp_ivl_25282;
  new_AGEMA_signal_4075 <= tmp_ivl_25289(1);
  n3920 <= tmp_ivl_25289(0);
  tmp_ivl_25289 <= LPM_d0_ivl_25293(0 + 1 downto 0);
  tmp_ivl_25294 <= new_AGEMA_signal_4075 & n3920;
  LPM_q_ivl_25297 <= tmp_ivl_25299 & tmp_ivl_25294;
  tmp_ivl_25301 <= new_AGEMA_signal_3763 & n3919;
  LPM_q_ivl_25304 <= tmp_ivl_25306 & tmp_ivl_25301;
  tmp_ivl_25308 <= tmp_ivl_25312(1);
  tmp_ivl_25310 <= tmp_ivl_25312(0);
  tmp_ivl_25312 <= LPM_d0_ivl_25316(0 + 1 downto 0);
  tmp_ivl_25317 <= new_AGEMA_signal_3648 & n3922;
  LPM_q_ivl_25320 <= tmp_ivl_25322 & tmp_ivl_25317;
  tmp_ivl_25324 <= new_AGEMA_signal_3707 & n3921;
  LPM_q_ivl_25327 <= tmp_ivl_25329 & tmp_ivl_25324;
  new_AGEMA_signal_4076 <= tmp_ivl_25331(1);
  n3924 <= tmp_ivl_25331(0);
  tmp_ivl_25331 <= LPM_d0_ivl_25335(0 + 1 downto 0);
  tmp_ivl_25337 <= state_in_s1(268);
  tmp_ivl_25339 <= state_in_s0(268);
  tmp_ivl_25340 <= tmp_ivl_25337 & tmp_ivl_25339;
  LPM_q_ivl_25343 <= tmp_ivl_25345 & tmp_ivl_25340;
  tmp_ivl_25347 <= new_AGEMA_signal_3453 & n3923;
  LPM_q_ivl_25350 <= tmp_ivl_25352 & tmp_ivl_25347;
  new_AGEMA_signal_3764 <= tmp_ivl_25354(1);
  n3930 <= tmp_ivl_25354(0);
  tmp_ivl_25354 <= LPM_d0_ivl_25358(0 + 1 downto 0);
  tmp_ivl_25359 <= new_AGEMA_signal_4076 & n3924;
  LPM_q_ivl_25362 <= tmp_ivl_25364 & tmp_ivl_25359;
  tmp_ivl_25366 <= new_AGEMA_signal_3764 & n3930;
  LPM_q_ivl_25369 <= tmp_ivl_25371 & tmp_ivl_25366;
  tmp_ivl_25373 <= tmp_ivl_25377(1);
  tmp_ivl_25375 <= tmp_ivl_25377(0);
  tmp_ivl_25377 <= LPM_d0_ivl_25381(0 + 1 downto 0);
  tmp_ivl_25382 <= new_AGEMA_signal_3585 & n3926;
  LPM_q_ivl_25385 <= tmp_ivl_25387 & tmp_ivl_25382;
  tmp_ivl_25389 <= new_AGEMA_signal_3598 & n3925;
  LPM_q_ivl_25392 <= tmp_ivl_25394 & tmp_ivl_25389;
  new_AGEMA_signal_4077 <= tmp_ivl_25396(1);
  n3927 <= tmp_ivl_25396(0);
  tmp_ivl_25396 <= LPM_d0_ivl_25400(0 + 1 downto 0);
  tmp_ivl_25401 <= new_AGEMA_signal_4077 & n3927;
  LPM_q_ivl_25404 <= tmp_ivl_25406 & tmp_ivl_25401;
  tmp_ivl_25408 <= new_AGEMA_signal_3764 & n3930;
  LPM_q_ivl_25411 <= tmp_ivl_25413 & tmp_ivl_25408;
  tmp_ivl_25415 <= tmp_ivl_25419(1);
  tmp_ivl_25417 <= tmp_ivl_25419(0);
  tmp_ivl_25419 <= LPM_d0_ivl_25423(0 + 1 downto 0);
  tmp_ivl_25424 <= new_AGEMA_signal_3597 & n3929;
  LPM_q_ivl_25427 <= tmp_ivl_25429 & tmp_ivl_25424;
  tmp_ivl_25431 <= new_AGEMA_signal_3760 & n3928;
  LPM_q_ivl_25434 <= tmp_ivl_25436 & tmp_ivl_25431;
  new_AGEMA_signal_4078 <= tmp_ivl_25438(1);
  n3931 <= tmp_ivl_25438(0);
  tmp_ivl_25438 <= LPM_d0_ivl_25442(0 + 1 downto 0);
  tmp_ivl_25443 <= new_AGEMA_signal_4078 & n3931;
  LPM_q_ivl_25446 <= tmp_ivl_25448 & tmp_ivl_25443;
  tmp_ivl_25450 <= new_AGEMA_signal_3764 & n3930;
  LPM_q_ivl_25453 <= tmp_ivl_25455 & tmp_ivl_25450;
  tmp_ivl_25457 <= tmp_ivl_25461(1);
  tmp_ivl_25459 <= tmp_ivl_25461(0);
  tmp_ivl_25461 <= LPM_d0_ivl_25465(0 + 1 downto 0);
  tmp_ivl_25466 <= new_AGEMA_signal_2692 & n3291;
  LPM_q_ivl_25469 <= tmp_ivl_25471 & tmp_ivl_25466;
  tmp_ivl_25474 <= z2(9);
  tmp_ivl_25475 <= new_AGEMA_signal_3292 & tmp_ivl_25474;
  LPM_q_ivl_25478 <= tmp_ivl_25480 & tmp_ivl_25475;
  new_AGEMA_signal_3454 <= tmp_ivl_25482(1);
  n4213 <= tmp_ivl_25482(0);
  tmp_ivl_25482 <= LPM_d0_ivl_25486(0 + 1 downto 0);
  tmp_ivl_25488 <= z3(9);
  tmp_ivl_25489 <= new_AGEMA_signal_3582 & tmp_ivl_25488;
  LPM_q_ivl_25492 <= tmp_ivl_25494 & tmp_ivl_25489;
  tmp_ivl_25497 <= state_in_s1(241);
  tmp_ivl_25499 <= state_in_s0(241);
  tmp_ivl_25500 <= tmp_ivl_25497 & tmp_ivl_25499;
  LPM_q_ivl_25503 <= tmp_ivl_25505 & tmp_ivl_25500;
  new_AGEMA_signal_3765 <= tmp_ivl_25507(1);
  n3932 <= tmp_ivl_25507(0);
  tmp_ivl_25507 <= LPM_d0_ivl_25511(0 + 1 downto 0);
  tmp_ivl_25512 <= new_AGEMA_signal_3454 & n4213;
  LPM_q_ivl_25515 <= tmp_ivl_25517 & tmp_ivl_25512;
  tmp_ivl_25519 <= new_AGEMA_signal_3765 & n3932;
  LPM_q_ivl_25522 <= tmp_ivl_25524 & tmp_ivl_25519;
  new_AGEMA_signal_4079 <= tmp_ivl_25526(1);
  n4072 <= tmp_ivl_25526(0);
  tmp_ivl_25526 <= LPM_d0_ivl_25530(0 + 1 downto 0);
  tmp_ivl_25531 <= new_AGEMA_signal_2695 & n3280;
  LPM_q_ivl_25534 <= tmp_ivl_25536 & tmp_ivl_25531;
  tmp_ivl_25539 <= z2(19);
  tmp_ivl_25540 <= new_AGEMA_signal_3282 & tmp_ivl_25539;
  LPM_q_ivl_25543 <= tmp_ivl_25545 & tmp_ivl_25540;
  new_AGEMA_signal_3455 <= tmp_ivl_25547(1);
  n4189 <= tmp_ivl_25547(0);
  tmp_ivl_25547 <= LPM_d0_ivl_25551(0 + 1 downto 0);
  tmp_ivl_25553 <= z3(19);
  tmp_ivl_25554 <= new_AGEMA_signal_3529 & tmp_ivl_25553;
  LPM_q_ivl_25557 <= tmp_ivl_25559 & tmp_ivl_25554;
  tmp_ivl_25562 <= state_in_s1(235);
  tmp_ivl_25564 <= state_in_s0(235);
  tmp_ivl_25565 <= tmp_ivl_25562 & tmp_ivl_25564;
  LPM_q_ivl_25568 <= tmp_ivl_25570 & tmp_ivl_25565;
  new_AGEMA_signal_3766 <= tmp_ivl_25572(1);
  n3933 <= tmp_ivl_25572(0);
  tmp_ivl_25572 <= LPM_d0_ivl_25576(0 + 1 downto 0);
  tmp_ivl_25577 <= new_AGEMA_signal_3455 & n4189;
  LPM_q_ivl_25580 <= tmp_ivl_25582 & tmp_ivl_25577;
  tmp_ivl_25584 <= new_AGEMA_signal_3766 & n3933;
  LPM_q_ivl_25587 <= tmp_ivl_25589 & tmp_ivl_25584;
  new_AGEMA_signal_4080 <= tmp_ivl_25591(1);
  n4076 <= tmp_ivl_25591(0);
  tmp_ivl_25591 <= LPM_d0_ivl_25595(0 + 1 downto 0);
  tmp_ivl_25596 <= new_AGEMA_signal_4079 & n4072;
  LPM_q_ivl_25599 <= tmp_ivl_25601 & tmp_ivl_25596;
  tmp_ivl_25603 <= new_AGEMA_signal_4080 & n4076;
  LPM_q_ivl_25606 <= tmp_ivl_25608 & tmp_ivl_25603;
  new_AGEMA_signal_4383 <= tmp_ivl_25610(1);
  n3935 <= tmp_ivl_25610(0);
  tmp_ivl_25610 <= LPM_d0_ivl_25614(0 + 1 downto 0);
  tmp_ivl_25615 <= new_AGEMA_signal_2698 & n3273;
  LPM_q_ivl_25618 <= tmp_ivl_25620 & tmp_ivl_25615;
  tmp_ivl_25623 <= z2(26);
  tmp_ivl_25624 <= new_AGEMA_signal_3293 & tmp_ivl_25623;
  LPM_q_ivl_25627 <= tmp_ivl_25629 & tmp_ivl_25624;
  new_AGEMA_signal_3456 <= tmp_ivl_25631(1);
  n4174 <= tmp_ivl_25631(0);
  tmp_ivl_25631 <= LPM_d0_ivl_25635(0 + 1 downto 0);
  tmp_ivl_25637 <= z3(26);
  tmp_ivl_25638 <= new_AGEMA_signal_3537 & tmp_ivl_25637;
  LPM_q_ivl_25641 <= tmp_ivl_25643 & tmp_ivl_25638;
  tmp_ivl_25646 <= state_in_s1(226);
  tmp_ivl_25648 <= state_in_s0(226);
  tmp_ivl_25649 <= tmp_ivl_25646 & tmp_ivl_25648;
  LPM_q_ivl_25652 <= tmp_ivl_25654 & tmp_ivl_25649;
  new_AGEMA_signal_3767 <= tmp_ivl_25656(1);
  n3934 <= tmp_ivl_25656(0);
  tmp_ivl_25656 <= LPM_d0_ivl_25660(0 + 1 downto 0);
  tmp_ivl_25661 <= new_AGEMA_signal_3456 & n4174;
  LPM_q_ivl_25664 <= tmp_ivl_25666 & tmp_ivl_25661;
  tmp_ivl_25668 <= new_AGEMA_signal_3767 & n3934;
  LPM_q_ivl_25671 <= tmp_ivl_25673 & tmp_ivl_25668;
  new_AGEMA_signal_4081 <= tmp_ivl_25675(1);
  n3984 <= tmp_ivl_25675(0);
  tmp_ivl_25675 <= LPM_d0_ivl_25679(0 + 1 downto 0);
  tmp_ivl_25680 <= new_AGEMA_signal_4383 & n3935;
  LPM_q_ivl_25683 <= tmp_ivl_25685 & tmp_ivl_25680;
  tmp_ivl_25687 <= new_AGEMA_signal_4081 & n3984;
  LPM_q_ivl_25690 <= tmp_ivl_25692 & tmp_ivl_25687;
  tmp_ivl_25694 <= tmp_ivl_25698(1);
  tmp_ivl_25696 <= tmp_ivl_25698(0);
  tmp_ivl_25698 <= LPM_d0_ivl_25702(0 + 1 downto 0);
  tmp_ivl_25703 <= new_AGEMA_signal_2701 & n3279;
  LPM_q_ivl_25706 <= tmp_ivl_25708 & tmp_ivl_25703;
  tmp_ivl_25711 <= z2(20);
  tmp_ivl_25712 <= new_AGEMA_signal_3279 & tmp_ivl_25711;
  LPM_q_ivl_25715 <= tmp_ivl_25717 & tmp_ivl_25712;
  new_AGEMA_signal_3457 <= tmp_ivl_25719(1);
  n4186 <= tmp_ivl_25719(0);
  tmp_ivl_25719 <= LPM_d0_ivl_25723(0 + 1 downto 0);
  tmp_ivl_25725 <= z3(20);
  tmp_ivl_25726 <= new_AGEMA_signal_3531 & tmp_ivl_25725;
  LPM_q_ivl_25729 <= tmp_ivl_25731 & tmp_ivl_25726;
  tmp_ivl_25734 <= state_in_s1(236);
  tmp_ivl_25736 <= state_in_s0(236);
  tmp_ivl_25737 <= tmp_ivl_25734 & tmp_ivl_25736;
  LPM_q_ivl_25740 <= tmp_ivl_25742 & tmp_ivl_25737;
  new_AGEMA_signal_3768 <= tmp_ivl_25744(1);
  n3936 <= tmp_ivl_25744(0);
  tmp_ivl_25744 <= LPM_d0_ivl_25748(0 + 1 downto 0);
  tmp_ivl_25749 <= new_AGEMA_signal_3457 & n4186;
  LPM_q_ivl_25752 <= tmp_ivl_25754 & tmp_ivl_25749;
  tmp_ivl_25756 <= new_AGEMA_signal_3768 & n3936;
  LPM_q_ivl_25759 <= tmp_ivl_25761 & tmp_ivl_25756;
  new_AGEMA_signal_4082 <= tmp_ivl_25763(1);
  n4264 <= tmp_ivl_25763(0);
  tmp_ivl_25763 <= LPM_d0_ivl_25767(0 + 1 downto 0);
  tmp_ivl_25768 <= new_AGEMA_signal_2704 & n3290;
  LPM_q_ivl_25771 <= tmp_ivl_25773 & tmp_ivl_25768;
  tmp_ivl_25776 <= z2(10);
  tmp_ivl_25777 <= new_AGEMA_signal_3285 & tmp_ivl_25776;
  LPM_q_ivl_25780 <= tmp_ivl_25782 & tmp_ivl_25777;
  new_AGEMA_signal_3458 <= tmp_ivl_25784(1);
  n4212 <= tmp_ivl_25784(0);
  tmp_ivl_25784 <= LPM_d0_ivl_25788(0 + 1 downto 0);
  tmp_ivl_25790 <= z3(10);
  tmp_ivl_25791 <= new_AGEMA_signal_3520 & tmp_ivl_25790;
  LPM_q_ivl_25794 <= tmp_ivl_25796 & tmp_ivl_25791;
  tmp_ivl_25799 <= state_in_s1(242);
  tmp_ivl_25801 <= state_in_s0(242);
  tmp_ivl_25802 <= tmp_ivl_25799 & tmp_ivl_25801;
  LPM_q_ivl_25805 <= tmp_ivl_25807 & tmp_ivl_25802;
  new_AGEMA_signal_3769 <= tmp_ivl_25809(1);
  n3937 <= tmp_ivl_25809(0);
  tmp_ivl_25809 <= LPM_d0_ivl_25813(0 + 1 downto 0);
  tmp_ivl_25814 <= new_AGEMA_signal_3458 & n4212;
  LPM_q_ivl_25817 <= tmp_ivl_25819 & tmp_ivl_25814;
  tmp_ivl_25821 <= new_AGEMA_signal_3769 & n3937;
  LPM_q_ivl_25824 <= tmp_ivl_25826 & tmp_ivl_25821;
  new_AGEMA_signal_4083 <= tmp_ivl_25828(1);
  n4269 <= tmp_ivl_25828(0);
  tmp_ivl_25828 <= LPM_d0_ivl_25832(0 + 1 downto 0);
  tmp_ivl_25833 <= new_AGEMA_signal_4082 & n4264;
  LPM_q_ivl_25836 <= tmp_ivl_25838 & tmp_ivl_25833;
  tmp_ivl_25840 <= new_AGEMA_signal_4083 & n4269;
  LPM_q_ivl_25843 <= tmp_ivl_25845 & tmp_ivl_25840;
  new_AGEMA_signal_4384 <= tmp_ivl_25847(1);
  n3939 <= tmp_ivl_25847(0);
  tmp_ivl_25847 <= LPM_d0_ivl_25851(0 + 1 downto 0);
  tmp_ivl_25852 <= new_AGEMA_signal_2707 & n3272;
  LPM_q_ivl_25855 <= tmp_ivl_25857 & tmp_ivl_25852;
  tmp_ivl_25860 <= z2(27);
  tmp_ivl_25861 <= new_AGEMA_signal_3291 & tmp_ivl_25860;
  LPM_q_ivl_25864 <= tmp_ivl_25866 & tmp_ivl_25861;
  new_AGEMA_signal_3459 <= tmp_ivl_25868(1);
  n4172 <= tmp_ivl_25868(0);
  tmp_ivl_25868 <= LPM_d0_ivl_25872(0 + 1 downto 0);
  tmp_ivl_25874 <= z3(27);
  tmp_ivl_25875 <= new_AGEMA_signal_3538 & tmp_ivl_25874;
  LPM_q_ivl_25878 <= tmp_ivl_25880 & tmp_ivl_25875;
  tmp_ivl_25883 <= state_in_s1(227);
  tmp_ivl_25885 <= state_in_s0(227);
  tmp_ivl_25886 <= tmp_ivl_25883 & tmp_ivl_25885;
  LPM_q_ivl_25889 <= tmp_ivl_25891 & tmp_ivl_25886;
  new_AGEMA_signal_3770 <= tmp_ivl_25893(1);
  n3938 <= tmp_ivl_25893(0);
  tmp_ivl_25893 <= LPM_d0_ivl_25897(0 + 1 downto 0);
  tmp_ivl_25898 <= new_AGEMA_signal_3459 & n4172;
  LPM_q_ivl_25901 <= tmp_ivl_25903 & tmp_ivl_25898;
  tmp_ivl_25905 <= new_AGEMA_signal_3770 & n3938;
  LPM_q_ivl_25908 <= tmp_ivl_25910 & tmp_ivl_25905;
  new_AGEMA_signal_4084 <= tmp_ivl_25912(1);
  n3987 <= tmp_ivl_25912(0);
  tmp_ivl_25912 <= LPM_d0_ivl_25916(0 + 1 downto 0);
  tmp_ivl_25917 <= new_AGEMA_signal_4384 & n3939;
  LPM_q_ivl_25920 <= tmp_ivl_25922 & tmp_ivl_25917;
  tmp_ivl_25924 <= new_AGEMA_signal_4084 & n3987;
  LPM_q_ivl_25927 <= tmp_ivl_25929 & tmp_ivl_25924;
  tmp_ivl_25931 <= tmp_ivl_25935(1);
  tmp_ivl_25933 <= tmp_ivl_25935(0);
  tmp_ivl_25935 <= LPM_d0_ivl_25939(0 + 1 downto 0);
  tmp_ivl_25940 <= new_AGEMA_signal_2709 & n3289;
  LPM_q_ivl_25943 <= tmp_ivl_25945 & tmp_ivl_25940;
  tmp_ivl_25948 <= z2(11);
  tmp_ivl_25949 <= new_AGEMA_signal_3283 & tmp_ivl_25948;
  LPM_q_ivl_25952 <= tmp_ivl_25954 & tmp_ivl_25949;
  new_AGEMA_signal_3460 <= tmp_ivl_25956(1);
  n4204 <= tmp_ivl_25956(0);
  tmp_ivl_25956 <= LPM_d0_ivl_25960(0 + 1 downto 0);
  tmp_ivl_25962 <= z3(11);
  tmp_ivl_25963 <= new_AGEMA_signal_3521 & tmp_ivl_25962;
  LPM_q_ivl_25966 <= tmp_ivl_25968 & tmp_ivl_25963;
  tmp_ivl_25971 <= state_in_s1(243);
  tmp_ivl_25973 <= state_in_s0(243);
  tmp_ivl_25974 <= tmp_ivl_25971 & tmp_ivl_25973;
  LPM_q_ivl_25977 <= tmp_ivl_25979 & tmp_ivl_25974;
  new_AGEMA_signal_3771 <= tmp_ivl_25981(1);
  n3940 <= tmp_ivl_25981(0);
  tmp_ivl_25981 <= LPM_d0_ivl_25985(0 + 1 downto 0);
  tmp_ivl_25986 <= new_AGEMA_signal_3460 & n4204;
  LPM_q_ivl_25989 <= tmp_ivl_25991 & tmp_ivl_25986;
  tmp_ivl_25993 <= new_AGEMA_signal_3771 & n3940;
  LPM_q_ivl_25996 <= tmp_ivl_25998 & tmp_ivl_25993;
  new_AGEMA_signal_4085 <= tmp_ivl_26000(1);
  n4258 <= tmp_ivl_26000(0);
  tmp_ivl_26000 <= LPM_d0_ivl_26004(0 + 1 downto 0);
  tmp_ivl_26005 <= new_AGEMA_signal_2712 & n3278;
  LPM_q_ivl_26008 <= tmp_ivl_26010 & tmp_ivl_26005;
  tmp_ivl_26013 <= z2(21);
  tmp_ivl_26014 <= new_AGEMA_signal_3278 & tmp_ivl_26013;
  LPM_q_ivl_26017 <= tmp_ivl_26019 & tmp_ivl_26014;
  new_AGEMA_signal_3461 <= tmp_ivl_26021(1);
  n4184 <= tmp_ivl_26021(0);
  tmp_ivl_26021 <= LPM_d0_ivl_26025(0 + 1 downto 0);
  tmp_ivl_26027 <= z3(21);
  tmp_ivl_26028 <= new_AGEMA_signal_3532 & tmp_ivl_26027;
  LPM_q_ivl_26031 <= tmp_ivl_26033 & tmp_ivl_26028;
  tmp_ivl_26036 <= state_in_s1(237);
  tmp_ivl_26038 <= state_in_s0(237);
  tmp_ivl_26039 <= tmp_ivl_26036 & tmp_ivl_26038;
  LPM_q_ivl_26042 <= tmp_ivl_26044 & tmp_ivl_26039;
  new_AGEMA_signal_3772 <= tmp_ivl_26046(1);
  n3941 <= tmp_ivl_26046(0);
  tmp_ivl_26046 <= LPM_d0_ivl_26050(0 + 1 downto 0);
  tmp_ivl_26051 <= new_AGEMA_signal_3461 & n4184;
  LPM_q_ivl_26054 <= tmp_ivl_26056 & tmp_ivl_26051;
  tmp_ivl_26058 <= new_AGEMA_signal_3772 & n3941;
  LPM_q_ivl_26061 <= tmp_ivl_26063 & tmp_ivl_26058;
  new_AGEMA_signal_4086 <= tmp_ivl_26065(1);
  n4254 <= tmp_ivl_26065(0);
  tmp_ivl_26065 <= LPM_d0_ivl_26069(0 + 1 downto 0);
  tmp_ivl_26070 <= new_AGEMA_signal_2714 & n3271;
  LPM_q_ivl_26073 <= tmp_ivl_26075 & tmp_ivl_26070;
  tmp_ivl_26078 <= z2(28);
  tmp_ivl_26079 <= new_AGEMA_signal_3290 & tmp_ivl_26078;
  LPM_q_ivl_26082 <= tmp_ivl_26084 & tmp_ivl_26079;
  new_AGEMA_signal_3462 <= tmp_ivl_26086(1);
  n4170 <= tmp_ivl_26086(0);
  tmp_ivl_26086 <= LPM_d0_ivl_26090(0 + 1 downto 0);
  tmp_ivl_26092 <= z3(28);
  tmp_ivl_26093 <= new_AGEMA_signal_3539 & tmp_ivl_26092;
  LPM_q_ivl_26096 <= tmp_ivl_26098 & tmp_ivl_26093;
  tmp_ivl_26101 <= state_in_s1(228);
  tmp_ivl_26103 <= state_in_s0(228);
  tmp_ivl_26104 <= tmp_ivl_26101 & tmp_ivl_26103;
  LPM_q_ivl_26107 <= tmp_ivl_26109 & tmp_ivl_26104;
  new_AGEMA_signal_3773 <= tmp_ivl_26111(1);
  n3942 <= tmp_ivl_26111(0);
  tmp_ivl_26111 <= LPM_d0_ivl_26115(0 + 1 downto 0);
  tmp_ivl_26116 <= new_AGEMA_signal_3462 & n4170;
  LPM_q_ivl_26119 <= tmp_ivl_26121 & tmp_ivl_26116;
  tmp_ivl_26123 <= new_AGEMA_signal_3773 & n3942;
  LPM_q_ivl_26126 <= tmp_ivl_26128 & tmp_ivl_26123;
  new_AGEMA_signal_4087 <= tmp_ivl_26130(1);
  n3989 <= tmp_ivl_26130(0);
  tmp_ivl_26130 <= LPM_d0_ivl_26134(0 + 1 downto 0);
  tmp_ivl_26135 <= new_AGEMA_signal_4086 & n4254;
  LPM_q_ivl_26138 <= tmp_ivl_26140 & tmp_ivl_26135;
  tmp_ivl_26142 <= new_AGEMA_signal_4087 & n3989;
  LPM_q_ivl_26145 <= tmp_ivl_26147 & tmp_ivl_26142;
  new_AGEMA_signal_4385 <= tmp_ivl_26149(1);
  n3943 <= tmp_ivl_26149(0);
  tmp_ivl_26149 <= LPM_d0_ivl_26153(0 + 1 downto 0);
  tmp_ivl_26154 <= new_AGEMA_signal_4085 & n4258;
  LPM_q_ivl_26157 <= tmp_ivl_26159 & tmp_ivl_26154;
  tmp_ivl_26161 <= new_AGEMA_signal_4385 & n3943;
  LPM_q_ivl_26164 <= tmp_ivl_26166 & tmp_ivl_26161;
  tmp_ivl_26168 <= tmp_ivl_26172(1);
  tmp_ivl_26170 <= tmp_ivl_26172(0);
  tmp_ivl_26172 <= LPM_d0_ivl_26176(0 + 1 downto 0);
  tmp_ivl_26177 <= new_AGEMA_signal_2717 & n3288;
  LPM_q_ivl_26180 <= tmp_ivl_26182 & tmp_ivl_26177;
  tmp_ivl_26185 <= z2(12);
  tmp_ivl_26186 <= new_AGEMA_signal_3281 & tmp_ivl_26185;
  LPM_q_ivl_26189 <= tmp_ivl_26191 & tmp_ivl_26186;
  new_AGEMA_signal_3463 <= tmp_ivl_26193(1);
  n4192 <= tmp_ivl_26193(0);
  tmp_ivl_26193 <= LPM_d0_ivl_26197(0 + 1 downto 0);
  tmp_ivl_26199 <= z3(12);
  tmp_ivl_26200 <= new_AGEMA_signal_3522 & tmp_ivl_26199;
  LPM_q_ivl_26203 <= tmp_ivl_26205 & tmp_ivl_26200;
  tmp_ivl_26208 <= state_in_s1(244);
  tmp_ivl_26210 <= state_in_s0(244);
  tmp_ivl_26211 <= tmp_ivl_26208 & tmp_ivl_26210;
  LPM_q_ivl_26214 <= tmp_ivl_26216 & tmp_ivl_26211;
  new_AGEMA_signal_3774 <= tmp_ivl_26218(1);
  n3944 <= tmp_ivl_26218(0);
  tmp_ivl_26218 <= LPM_d0_ivl_26222(0 + 1 downto 0);
  tmp_ivl_26223 <= new_AGEMA_signal_3463 & n4192;
  LPM_q_ivl_26226 <= tmp_ivl_26228 & tmp_ivl_26223;
  tmp_ivl_26230 <= new_AGEMA_signal_3774 & n3944;
  LPM_q_ivl_26233 <= tmp_ivl_26235 & tmp_ivl_26230;
  new_AGEMA_signal_4088 <= tmp_ivl_26237(1);
  n4245 <= tmp_ivl_26237(0);
  tmp_ivl_26237 <= LPM_d0_ivl_26241(0 + 1 downto 0);
  tmp_ivl_26242 <= new_AGEMA_signal_2719 & n3277;
  LPM_q_ivl_26245 <= tmp_ivl_26247 & tmp_ivl_26242;
  tmp_ivl_26250 <= z2(22);
  tmp_ivl_26251 <= new_AGEMA_signal_3275 & tmp_ivl_26250;
  LPM_q_ivl_26254 <= tmp_ivl_26256 & tmp_ivl_26251;
  new_AGEMA_signal_3464 <= tmp_ivl_26258(1);
  n4183 <= tmp_ivl_26258(0);
  tmp_ivl_26258 <= LPM_d0_ivl_26262(0 + 1 downto 0);
  tmp_ivl_26264 <= z3(22);
  tmp_ivl_26265 <= new_AGEMA_signal_3533 & tmp_ivl_26264;
  LPM_q_ivl_26268 <= tmp_ivl_26270 & tmp_ivl_26265;
  tmp_ivl_26273 <= state_in_s1(238);
  tmp_ivl_26275 <= state_in_s0(238);
  tmp_ivl_26276 <= tmp_ivl_26273 & tmp_ivl_26275;
  LPM_q_ivl_26279 <= tmp_ivl_26281 & tmp_ivl_26276;
  new_AGEMA_signal_3775 <= tmp_ivl_26283(1);
  n3945 <= tmp_ivl_26283(0);
  tmp_ivl_26283 <= LPM_d0_ivl_26287(0 + 1 downto 0);
  tmp_ivl_26288 <= new_AGEMA_signal_3464 & n4183;
  LPM_q_ivl_26291 <= tmp_ivl_26293 & tmp_ivl_26288;
  tmp_ivl_26295 <= new_AGEMA_signal_3775 & n3945;
  LPM_q_ivl_26298 <= tmp_ivl_26300 & tmp_ivl_26295;
  new_AGEMA_signal_4089 <= tmp_ivl_26302(1);
  n4241 <= tmp_ivl_26302(0);
  tmp_ivl_26302 <= LPM_d0_ivl_26306(0 + 1 downto 0);
  tmp_ivl_26307 <= new_AGEMA_signal_2721 & n3270;
  LPM_q_ivl_26310 <= tmp_ivl_26312 & tmp_ivl_26307;
  tmp_ivl_26315 <= z2(29);
  tmp_ivl_26316 <= new_AGEMA_signal_3289 & tmp_ivl_26315;
  LPM_q_ivl_26319 <= tmp_ivl_26321 & tmp_ivl_26316;
  new_AGEMA_signal_3465 <= tmp_ivl_26323(1);
  n4169 <= tmp_ivl_26323(0);
  tmp_ivl_26323 <= LPM_d0_ivl_26327(0 + 1 downto 0);
  tmp_ivl_26329 <= z3(29);
  tmp_ivl_26330 <= new_AGEMA_signal_3540 & tmp_ivl_26329;
  LPM_q_ivl_26333 <= tmp_ivl_26335 & tmp_ivl_26330;
  tmp_ivl_26338 <= state_in_s1(229);
  tmp_ivl_26340 <= state_in_s0(229);
  tmp_ivl_26341 <= tmp_ivl_26338 & tmp_ivl_26340;
  LPM_q_ivl_26344 <= tmp_ivl_26346 & tmp_ivl_26341;
  new_AGEMA_signal_3776 <= tmp_ivl_26348(1);
  n3946 <= tmp_ivl_26348(0);
  tmp_ivl_26348 <= LPM_d0_ivl_26352(0 + 1 downto 0);
  tmp_ivl_26353 <= new_AGEMA_signal_3465 & n4169;
  LPM_q_ivl_26356 <= tmp_ivl_26358 & tmp_ivl_26353;
  tmp_ivl_26360 <= new_AGEMA_signal_3776 & n3946;
  LPM_q_ivl_26363 <= tmp_ivl_26365 & tmp_ivl_26360;
  new_AGEMA_signal_4090 <= tmp_ivl_26367(1);
  n3992 <= tmp_ivl_26367(0);
  tmp_ivl_26367 <= LPM_d0_ivl_26371(0 + 1 downto 0);
  tmp_ivl_26372 <= new_AGEMA_signal_4089 & n4241;
  LPM_q_ivl_26375 <= tmp_ivl_26377 & tmp_ivl_26372;
  tmp_ivl_26379 <= new_AGEMA_signal_4090 & n3992;
  LPM_q_ivl_26382 <= tmp_ivl_26384 & tmp_ivl_26379;
  new_AGEMA_signal_4386 <= tmp_ivl_26386(1);
  n3947 <= tmp_ivl_26386(0);
  tmp_ivl_26386 <= LPM_d0_ivl_26390(0 + 1 downto 0);
  tmp_ivl_26391 <= new_AGEMA_signal_4088 & n4245;
  LPM_q_ivl_26394 <= tmp_ivl_26396 & tmp_ivl_26391;
  tmp_ivl_26398 <= new_AGEMA_signal_4386 & n3947;
  LPM_q_ivl_26401 <= tmp_ivl_26403 & tmp_ivl_26398;
  tmp_ivl_26405 <= tmp_ivl_26409(1);
  tmp_ivl_26407 <= tmp_ivl_26409(0);
  tmp_ivl_26409 <= LPM_d0_ivl_26413(0 + 1 downto 0);
  tmp_ivl_26414 <= new_AGEMA_signal_2724 & n3276;
  LPM_q_ivl_26417 <= tmp_ivl_26419 & tmp_ivl_26414;
  tmp_ivl_26422 <= z2(23);
  tmp_ivl_26423 <= new_AGEMA_signal_3273 & tmp_ivl_26422;
  LPM_q_ivl_26426 <= tmp_ivl_26428 & tmp_ivl_26423;
  new_AGEMA_signal_3466 <= tmp_ivl_26430(1);
  n4180 <= tmp_ivl_26430(0);
  tmp_ivl_26430 <= LPM_d0_ivl_26434(0 + 1 downto 0);
  tmp_ivl_26436 <= z3(23);
  tmp_ivl_26437 <= new_AGEMA_signal_3534 & tmp_ivl_26436;
  LPM_q_ivl_26440 <= tmp_ivl_26442 & tmp_ivl_26437;
  tmp_ivl_26445 <= state_in_s1(239);
  tmp_ivl_26447 <= state_in_s0(239);
  tmp_ivl_26448 <= tmp_ivl_26445 & tmp_ivl_26447;
  LPM_q_ivl_26451 <= tmp_ivl_26453 & tmp_ivl_26448;
  new_AGEMA_signal_3777 <= tmp_ivl_26455(1);
  n3948 <= tmp_ivl_26455(0);
  tmp_ivl_26455 <= LPM_d0_ivl_26459(0 + 1 downto 0);
  tmp_ivl_26460 <= new_AGEMA_signal_3466 & n4180;
  LPM_q_ivl_26463 <= tmp_ivl_26465 & tmp_ivl_26460;
  tmp_ivl_26467 <= new_AGEMA_signal_3777 & n3948;
  LPM_q_ivl_26470 <= tmp_ivl_26472 & tmp_ivl_26467;
  new_AGEMA_signal_4091 <= tmp_ivl_26474(1);
  n4230 <= tmp_ivl_26474(0);
  tmp_ivl_26474 <= LPM_d0_ivl_26478(0 + 1 downto 0);
  tmp_ivl_26479 <= new_AGEMA_signal_2727 & n3286;
  LPM_q_ivl_26482 <= tmp_ivl_26484 & tmp_ivl_26479;
  tmp_ivl_26487 <= z2(13);
  tmp_ivl_26488 <= new_AGEMA_signal_3280 & tmp_ivl_26487;
  LPM_q_ivl_26491 <= tmp_ivl_26493 & tmp_ivl_26488;
  new_AGEMA_signal_3467 <= tmp_ivl_26495(1);
  n4201 <= tmp_ivl_26495(0);
  tmp_ivl_26495 <= LPM_d0_ivl_26499(0 + 1 downto 0);
  tmp_ivl_26501 <= z3(13);
  tmp_ivl_26502 <= new_AGEMA_signal_3523 & tmp_ivl_26501;
  LPM_q_ivl_26505 <= tmp_ivl_26507 & tmp_ivl_26502;
  tmp_ivl_26510 <= state_in_s1(245);
  tmp_ivl_26512 <= state_in_s0(245);
  tmp_ivl_26513 <= tmp_ivl_26510 & tmp_ivl_26512;
  LPM_q_ivl_26516 <= tmp_ivl_26518 & tmp_ivl_26513;
  new_AGEMA_signal_3778 <= tmp_ivl_26520(1);
  n3949 <= tmp_ivl_26520(0);
  tmp_ivl_26520 <= LPM_d0_ivl_26524(0 + 1 downto 0);
  tmp_ivl_26525 <= new_AGEMA_signal_3467 & n4201;
  LPM_q_ivl_26528 <= tmp_ivl_26530 & tmp_ivl_26525;
  tmp_ivl_26532 <= new_AGEMA_signal_3778 & n3949;
  LPM_q_ivl_26535 <= tmp_ivl_26537 & tmp_ivl_26532;
  new_AGEMA_signal_4092 <= tmp_ivl_26539(1);
  n4263 <= tmp_ivl_26539(0);
  tmp_ivl_26539 <= LPM_d0_ivl_26543(0 + 1 downto 0);
  tmp_ivl_26544 <= new_AGEMA_signal_4091 & n4230;
  LPM_q_ivl_26547 <= tmp_ivl_26549 & tmp_ivl_26544;
  tmp_ivl_26551 <= new_AGEMA_signal_4092 & n4263;
  LPM_q_ivl_26554 <= tmp_ivl_26556 & tmp_ivl_26551;
  new_AGEMA_signal_4387 <= tmp_ivl_26558(1);
  n3951 <= tmp_ivl_26558(0);
  tmp_ivl_26558 <= LPM_d0_ivl_26562(0 + 1 downto 0);
  tmp_ivl_26563 <= new_AGEMA_signal_2730 & n3269;
  LPM_q_ivl_26566 <= tmp_ivl_26568 & tmp_ivl_26563;
  tmp_ivl_26571 <= z2(30);
  tmp_ivl_26572 <= new_AGEMA_signal_3288 & tmp_ivl_26571;
  LPM_q_ivl_26575 <= tmp_ivl_26577 & tmp_ivl_26572;
  new_AGEMA_signal_3468 <= tmp_ivl_26579(1);
  n4166 <= tmp_ivl_26579(0);
  tmp_ivl_26579 <= LPM_d0_ivl_26583(0 + 1 downto 0);
  tmp_ivl_26585 <= z3(30);
  tmp_ivl_26586 <= new_AGEMA_signal_3542 & tmp_ivl_26585;
  LPM_q_ivl_26589 <= tmp_ivl_26591 & tmp_ivl_26586;
  tmp_ivl_26594 <= state_in_s1(230);
  tmp_ivl_26596 <= state_in_s0(230);
  tmp_ivl_26597 <= tmp_ivl_26594 & tmp_ivl_26596;
  LPM_q_ivl_26600 <= tmp_ivl_26602 & tmp_ivl_26597;
  new_AGEMA_signal_3779 <= tmp_ivl_26604(1);
  n3950 <= tmp_ivl_26604(0);
  tmp_ivl_26604 <= LPM_d0_ivl_26608(0 + 1 downto 0);
  tmp_ivl_26609 <= new_AGEMA_signal_3468 & n4166;
  LPM_q_ivl_26612 <= tmp_ivl_26614 & tmp_ivl_26609;
  tmp_ivl_26616 <= new_AGEMA_signal_3779 & n3950;
  LPM_q_ivl_26619 <= tmp_ivl_26621 & tmp_ivl_26616;
  new_AGEMA_signal_4093 <= tmp_ivl_26623(1);
  n3996 <= tmp_ivl_26623(0);
  tmp_ivl_26623 <= LPM_d0_ivl_26627(0 + 1 downto 0);
  tmp_ivl_26628 <= new_AGEMA_signal_4387 & n3951;
  LPM_q_ivl_26631 <= tmp_ivl_26633 & tmp_ivl_26628;
  tmp_ivl_26635 <= new_AGEMA_signal_4093 & n3996;
  LPM_q_ivl_26638 <= tmp_ivl_26640 & tmp_ivl_26635;
  tmp_ivl_26642 <= tmp_ivl_26646(1);
  tmp_ivl_26644 <= tmp_ivl_26646(0);
  tmp_ivl_26646 <= LPM_d0_ivl_26650(0 + 1 downto 0);
  tmp_ivl_26651 <= new_AGEMA_signal_2733 & n3285;
  LPM_q_ivl_26654 <= tmp_ivl_26656 & tmp_ivl_26651;
  tmp_ivl_26659 <= z2(14);
  tmp_ivl_26660 <= new_AGEMA_signal_3277 & tmp_ivl_26659;
  LPM_q_ivl_26663 <= tmp_ivl_26665 & tmp_ivl_26660;
  new_AGEMA_signal_3469 <= tmp_ivl_26667(1);
  n4199 <= tmp_ivl_26667(0);
  tmp_ivl_26667 <= LPM_d0_ivl_26671(0 + 1 downto 0);
  tmp_ivl_26673 <= z3(14);
  tmp_ivl_26674 <= new_AGEMA_signal_3524 & tmp_ivl_26673;
  LPM_q_ivl_26677 <= tmp_ivl_26679 & tmp_ivl_26674;
  tmp_ivl_26682 <= state_in_s1(246);
  tmp_ivl_26684 <= state_in_s0(246);
  tmp_ivl_26685 <= tmp_ivl_26682 & tmp_ivl_26684;
  LPM_q_ivl_26688 <= tmp_ivl_26690 & tmp_ivl_26685;
  new_AGEMA_signal_3780 <= tmp_ivl_26692(1);
  n3952 <= tmp_ivl_26692(0);
  tmp_ivl_26692 <= LPM_d0_ivl_26696(0 + 1 downto 0);
  tmp_ivl_26697 <= new_AGEMA_signal_3469 & n4199;
  LPM_q_ivl_26700 <= tmp_ivl_26702 & tmp_ivl_26697;
  tmp_ivl_26704 <= new_AGEMA_signal_3780 & n3952;
  LPM_q_ivl_26707 <= tmp_ivl_26709 & tmp_ivl_26704;
  new_AGEMA_signal_4094 <= tmp_ivl_26711(1);
  n4255 <= tmp_ivl_26711(0);
  tmp_ivl_26711 <= LPM_d0_ivl_26715(0 + 1 downto 0);
  tmp_ivl_26716 <= new_AGEMA_signal_2736 & n3275;
  LPM_q_ivl_26719 <= tmp_ivl_26721 & tmp_ivl_26716;
  tmp_ivl_26724 <= z2(24);
  tmp_ivl_26725 <= new_AGEMA_signal_3271 & tmp_ivl_26724;
  LPM_q_ivl_26728 <= tmp_ivl_26730 & tmp_ivl_26725;
  new_AGEMA_signal_3470 <= tmp_ivl_26732(1);
  n4178 <= tmp_ivl_26732(0);
  tmp_ivl_26732 <= LPM_d0_ivl_26736(0 + 1 downto 0);
  tmp_ivl_26738 <= z3(24);
  tmp_ivl_26739 <= new_AGEMA_signal_3535 & tmp_ivl_26738;
  LPM_q_ivl_26742 <= tmp_ivl_26744 & tmp_ivl_26739;
  tmp_ivl_26747 <= state_in_s1(224);
  tmp_ivl_26749 <= state_in_s0(224);
  tmp_ivl_26750 <= tmp_ivl_26747 & tmp_ivl_26749;
  LPM_q_ivl_26753 <= tmp_ivl_26755 & tmp_ivl_26750;
  new_AGEMA_signal_3781 <= tmp_ivl_26757(1);
  n3953 <= tmp_ivl_26757(0);
  tmp_ivl_26757 <= LPM_d0_ivl_26761(0 + 1 downto 0);
  tmp_ivl_26762 <= new_AGEMA_signal_3470 & n4178;
  LPM_q_ivl_26765 <= tmp_ivl_26767 & tmp_ivl_26762;
  tmp_ivl_26769 <= new_AGEMA_signal_3781 & n3953;
  LPM_q_ivl_26772 <= tmp_ivl_26774 & tmp_ivl_26769;
  new_AGEMA_signal_4095 <= tmp_ivl_26776(1);
  n4094 <= tmp_ivl_26776(0);
  tmp_ivl_26776 <= LPM_d0_ivl_26780(0 + 1 downto 0);
  tmp_ivl_26781 <= new_AGEMA_signal_4094 & n4255;
  LPM_q_ivl_26784 <= tmp_ivl_26786 & tmp_ivl_26781;
  tmp_ivl_26788 <= new_AGEMA_signal_4095 & n4094;
  LPM_q_ivl_26791 <= tmp_ivl_26793 & tmp_ivl_26788;
  new_AGEMA_signal_4388 <= tmp_ivl_26795(1);
  n3955 <= tmp_ivl_26795(0);
  tmp_ivl_26795 <= LPM_d0_ivl_26799(0 + 1 downto 0);
  tmp_ivl_26800 <= new_AGEMA_signal_2739 & n3268;
  LPM_q_ivl_26803 <= tmp_ivl_26805 & tmp_ivl_26800;
  tmp_ivl_26808 <= z2(31);
  tmp_ivl_26809 <= new_AGEMA_signal_3287 & tmp_ivl_26808;
  LPM_q_ivl_26812 <= tmp_ivl_26814 & tmp_ivl_26809;
  new_AGEMA_signal_3471 <= tmp_ivl_26816(1);
  n4164 <= tmp_ivl_26816(0);
  tmp_ivl_26816 <= LPM_d0_ivl_26820(0 + 1 downto 0);
  tmp_ivl_26822 <= z3(31);
  tmp_ivl_26823 <= new_AGEMA_signal_3543 & tmp_ivl_26822;
  LPM_q_ivl_26826 <= tmp_ivl_26828 & tmp_ivl_26823;
  tmp_ivl_26831 <= state_in_s1(231);
  tmp_ivl_26833 <= state_in_s0(231);
  tmp_ivl_26834 <= tmp_ivl_26831 & tmp_ivl_26833;
  LPM_q_ivl_26837 <= tmp_ivl_26839 & tmp_ivl_26834;
  new_AGEMA_signal_3782 <= tmp_ivl_26841(1);
  n3954 <= tmp_ivl_26841(0);
  tmp_ivl_26841 <= LPM_d0_ivl_26845(0 + 1 downto 0);
  tmp_ivl_26846 <= new_AGEMA_signal_3471 & n4164;
  LPM_q_ivl_26849 <= tmp_ivl_26851 & tmp_ivl_26846;
  tmp_ivl_26853 <= new_AGEMA_signal_3782 & n3954;
  LPM_q_ivl_26856 <= tmp_ivl_26858 & tmp_ivl_26853;
  new_AGEMA_signal_4096 <= tmp_ivl_26860(1);
  n3998 <= tmp_ivl_26860(0);
  tmp_ivl_26860 <= LPM_d0_ivl_26864(0 + 1 downto 0);
  tmp_ivl_26865 <= new_AGEMA_signal_4388 & n3955;
  LPM_q_ivl_26868 <= tmp_ivl_26870 & tmp_ivl_26865;
  tmp_ivl_26872 <= new_AGEMA_signal_4096 & n3998;
  LPM_q_ivl_26875 <= tmp_ivl_26877 & tmp_ivl_26872;
  tmp_ivl_26879 <= tmp_ivl_26883(1);
  tmp_ivl_26881 <= tmp_ivl_26883(0);
  tmp_ivl_26883 <= LPM_d0_ivl_26887(0 + 1 downto 0);
  tmp_ivl_26888 <= new_AGEMA_signal_2742 & n3284;
  LPM_q_ivl_26891 <= tmp_ivl_26893 & tmp_ivl_26888;
  tmp_ivl_26896 <= z2(15);
  tmp_ivl_26897 <= new_AGEMA_signal_3276 & tmp_ivl_26896;
  LPM_q_ivl_26900 <= tmp_ivl_26902 & tmp_ivl_26897;
  new_AGEMA_signal_3472 <= tmp_ivl_26904(1);
  n4198 <= tmp_ivl_26904(0);
  tmp_ivl_26904 <= LPM_d0_ivl_26908(0 + 1 downto 0);
  tmp_ivl_26910 <= z3(15);
  tmp_ivl_26911 <= new_AGEMA_signal_3525 & tmp_ivl_26910;
  LPM_q_ivl_26914 <= tmp_ivl_26916 & tmp_ivl_26911;
  tmp_ivl_26919 <= state_in_s1(247);
  tmp_ivl_26921 <= state_in_s0(247);
  tmp_ivl_26922 <= tmp_ivl_26919 & tmp_ivl_26921;
  LPM_q_ivl_26925 <= tmp_ivl_26927 & tmp_ivl_26922;
  new_AGEMA_signal_3783 <= tmp_ivl_26929(1);
  n3956 <= tmp_ivl_26929(0);
  tmp_ivl_26929 <= LPM_d0_ivl_26933(0 + 1 downto 0);
  tmp_ivl_26934 <= new_AGEMA_signal_3472 & n4198;
  LPM_q_ivl_26937 <= tmp_ivl_26939 & tmp_ivl_26934;
  tmp_ivl_26941 <= new_AGEMA_signal_3783 & n3956;
  LPM_q_ivl_26944 <= tmp_ivl_26946 & tmp_ivl_26941;
  new_AGEMA_signal_4097 <= tmp_ivl_26948(1);
  n4239 <= tmp_ivl_26948(0);
  tmp_ivl_26948 <= LPM_d0_ivl_26952(0 + 1 downto 0);
  tmp_ivl_26953 <= new_AGEMA_signal_2744 & n3274;
  LPM_q_ivl_26956 <= tmp_ivl_26958 & tmp_ivl_26953;
  tmp_ivl_26961 <= z2(25);
  tmp_ivl_26962 <= new_AGEMA_signal_3286 & tmp_ivl_26961;
  LPM_q_ivl_26965 <= tmp_ivl_26967 & tmp_ivl_26962;
  new_AGEMA_signal_3473 <= tmp_ivl_26969(1);
  n4177 <= tmp_ivl_26969(0);
  tmp_ivl_26969 <= LPM_d0_ivl_26973(0 + 1 downto 0);
  tmp_ivl_26975 <= z3(25);
  tmp_ivl_26976 <= new_AGEMA_signal_3536 & tmp_ivl_26975;
  LPM_q_ivl_26979 <= tmp_ivl_26981 & tmp_ivl_26976;
  tmp_ivl_26984 <= state_in_s1(225);
  tmp_ivl_26986 <= state_in_s0(225);
  tmp_ivl_26987 <= tmp_ivl_26984 & tmp_ivl_26986;
  LPM_q_ivl_26990 <= tmp_ivl_26992 & tmp_ivl_26987;
  new_AGEMA_signal_3784 <= tmp_ivl_26994(1);
  n3957 <= tmp_ivl_26994(0);
  tmp_ivl_26994 <= LPM_d0_ivl_26998(0 + 1 downto 0);
  tmp_ivl_26999 <= new_AGEMA_signal_3473 & n4177;
  LPM_q_ivl_27002 <= tmp_ivl_27004 & tmp_ivl_26999;
  tmp_ivl_27006 <= new_AGEMA_signal_3784 & n3957;
  LPM_q_ivl_27009 <= tmp_ivl_27011 & tmp_ivl_27006;
  new_AGEMA_signal_4098 <= tmp_ivl_27013(1);
  n4044 <= tmp_ivl_27013(0);
  tmp_ivl_27013 <= LPM_d0_ivl_27017(0 + 1 downto 0);
  tmp_ivl_27018 <= new_AGEMA_signal_2747 & n3267;
  LPM_q_ivl_27021 <= tmp_ivl_27023 & tmp_ivl_27018;
  tmp_ivl_27026 <= z2(32);
  tmp_ivl_27027 <= new_AGEMA_signal_3188 & tmp_ivl_27026;
  LPM_q_ivl_27030 <= tmp_ivl_27032 & tmp_ivl_27027;
  new_AGEMA_signal_3474 <= tmp_ivl_27034(1);
  n4163 <= tmp_ivl_27034(0);
  tmp_ivl_27034 <= LPM_d0_ivl_27038(0 + 1 downto 0);
  tmp_ivl_27040 <= z3(32);
  tmp_ivl_27041 <= new_AGEMA_signal_3544 & tmp_ivl_27040;
  LPM_q_ivl_27044 <= tmp_ivl_27046 & tmp_ivl_27041;
  tmp_ivl_27049 <= state_in_s1(216);
  tmp_ivl_27051 <= state_in_s0(216);
  tmp_ivl_27052 <= tmp_ivl_27049 & tmp_ivl_27051;
  LPM_q_ivl_27055 <= tmp_ivl_27057 & tmp_ivl_27052;
  new_AGEMA_signal_3785 <= tmp_ivl_27059(1);
  n3958 <= tmp_ivl_27059(0);
  tmp_ivl_27059 <= LPM_d0_ivl_27063(0 + 1 downto 0);
  tmp_ivl_27064 <= new_AGEMA_signal_3474 & n4163;
  LPM_q_ivl_27067 <= tmp_ivl_27069 & tmp_ivl_27064;
  tmp_ivl_27071 <= new_AGEMA_signal_3785 & n3958;
  LPM_q_ivl_27074 <= tmp_ivl_27076 & tmp_ivl_27071;
  new_AGEMA_signal_4099 <= tmp_ivl_27078(1);
  n4002 <= tmp_ivl_27078(0);
  tmp_ivl_27078 <= LPM_d0_ivl_27082(0 + 1 downto 0);
  tmp_ivl_27083 <= new_AGEMA_signal_4098 & n4044;
  LPM_q_ivl_27086 <= tmp_ivl_27088 & tmp_ivl_27083;
  tmp_ivl_27090 <= new_AGEMA_signal_4099 & n4002;
  LPM_q_ivl_27093 <= tmp_ivl_27095 & tmp_ivl_27090;
  new_AGEMA_signal_4389 <= tmp_ivl_27097(1);
  n3959 <= tmp_ivl_27097(0);
  tmp_ivl_27097 <= LPM_d0_ivl_27101(0 + 1 downto 0);
  tmp_ivl_27102 <= new_AGEMA_signal_4097 & n4239;
  LPM_q_ivl_27105 <= tmp_ivl_27107 & tmp_ivl_27102;
  tmp_ivl_27109 <= new_AGEMA_signal_4389 & n3959;
  LPM_q_ivl_27112 <= tmp_ivl_27114 & tmp_ivl_27109;
  tmp_ivl_27116 <= tmp_ivl_27120(1);
  tmp_ivl_27118 <= tmp_ivl_27120(0);
  tmp_ivl_27120 <= LPM_d0_ivl_27124(0 + 1 downto 0);
  tmp_ivl_27125 <= new_AGEMA_signal_2750 & n3283;
  LPM_q_ivl_27128 <= tmp_ivl_27130 & tmp_ivl_27125;
  tmp_ivl_27133 <= z2(16);
  tmp_ivl_27134 <= new_AGEMA_signal_3274 & tmp_ivl_27133;
  LPM_q_ivl_27137 <= tmp_ivl_27139 & tmp_ivl_27134;
  new_AGEMA_signal_3475 <= tmp_ivl_27141(1);
  n4195 <= tmp_ivl_27141(0);
  tmp_ivl_27141 <= LPM_d0_ivl_27145(0 + 1 downto 0);
  tmp_ivl_27147 <= z3(16);
  tmp_ivl_27148 <= new_AGEMA_signal_3526 & tmp_ivl_27147;
  LPM_q_ivl_27151 <= tmp_ivl_27153 & tmp_ivl_27148;
  tmp_ivl_27156 <= state_in_s1(232);
  tmp_ivl_27158 <= state_in_s0(232);
  tmp_ivl_27159 <= tmp_ivl_27156 & tmp_ivl_27158;
  LPM_q_ivl_27162 <= tmp_ivl_27164 & tmp_ivl_27159;
  new_AGEMA_signal_3786 <= tmp_ivl_27166(1);
  n3960 <= tmp_ivl_27166(0);
  tmp_ivl_27166 <= LPM_d0_ivl_27170(0 + 1 downto 0);
  tmp_ivl_27171 <= new_AGEMA_signal_3475 & n4195;
  LPM_q_ivl_27174 <= tmp_ivl_27176 & tmp_ivl_27171;
  tmp_ivl_27178 <= new_AGEMA_signal_3786 & n3960;
  LPM_q_ivl_27181 <= tmp_ivl_27183 & tmp_ivl_27178;
  new_AGEMA_signal_4100 <= tmp_ivl_27185(1);
  n4229 <= tmp_ivl_27185(0);
  tmp_ivl_27185 <= LPM_d0_ivl_27189(0 + 1 downto 0);
  tmp_ivl_27190 <= new_AGEMA_signal_4100 & n4229;
  LPM_q_ivl_27193 <= tmp_ivl_27195 & tmp_ivl_27190;
  tmp_ivl_27197 <= new_AGEMA_signal_4081 & n3984;
  LPM_q_ivl_27200 <= tmp_ivl_27202 & tmp_ivl_27197;
  new_AGEMA_signal_4390 <= tmp_ivl_27204(1);
  n3962 <= tmp_ivl_27204(0);
  tmp_ivl_27204 <= LPM_d0_ivl_27208(0 + 1 downto 0);
  tmp_ivl_27209 <= new_AGEMA_signal_2753 & n3266;
  LPM_q_ivl_27212 <= tmp_ivl_27214 & tmp_ivl_27209;
  tmp_ivl_27217 <= z2(33);
  tmp_ivl_27218 <= new_AGEMA_signal_3187 & tmp_ivl_27217;
  LPM_q_ivl_27221 <= tmp_ivl_27223 & tmp_ivl_27218;
  new_AGEMA_signal_3476 <= tmp_ivl_27225(1);
  n4161 <= tmp_ivl_27225(0);
  tmp_ivl_27225 <= LPM_d0_ivl_27229(0 + 1 downto 0);
  tmp_ivl_27231 <= z3(33);
  tmp_ivl_27232 <= new_AGEMA_signal_3545 & tmp_ivl_27231;
  LPM_q_ivl_27235 <= tmp_ivl_27237 & tmp_ivl_27232;
  tmp_ivl_27240 <= state_in_s1(217);
  tmp_ivl_27242 <= state_in_s0(217);
  tmp_ivl_27243 <= tmp_ivl_27240 & tmp_ivl_27242;
  LPM_q_ivl_27246 <= tmp_ivl_27248 & tmp_ivl_27243;
  new_AGEMA_signal_3787 <= tmp_ivl_27250(1);
  n3961 <= tmp_ivl_27250(0);
  tmp_ivl_27250 <= LPM_d0_ivl_27254(0 + 1 downto 0);
  tmp_ivl_27255 <= new_AGEMA_signal_3476 & n4161;
  LPM_q_ivl_27258 <= tmp_ivl_27260 & tmp_ivl_27255;
  tmp_ivl_27262 <= new_AGEMA_signal_3787 & n3961;
  LPM_q_ivl_27265 <= tmp_ivl_27267 & tmp_ivl_27262;
  new_AGEMA_signal_4101 <= tmp_ivl_27269(1);
  n4006 <= tmp_ivl_27269(0);
  tmp_ivl_27269 <= LPM_d0_ivl_27273(0 + 1 downto 0);
  tmp_ivl_27274 <= new_AGEMA_signal_4390 & n3962;
  LPM_q_ivl_27277 <= tmp_ivl_27279 & tmp_ivl_27274;
  tmp_ivl_27281 <= new_AGEMA_signal_4101 & n4006;
  LPM_q_ivl_27284 <= tmp_ivl_27286 & tmp_ivl_27281;
  tmp_ivl_27288 <= tmp_ivl_27292(1);
  tmp_ivl_27290 <= tmp_ivl_27292(0);
  tmp_ivl_27292 <= LPM_d0_ivl_27296(0 + 1 downto 0);
  tmp_ivl_27297 <= new_AGEMA_signal_2755 & n3282;
  LPM_q_ivl_27300 <= tmp_ivl_27302 & tmp_ivl_27297;
  tmp_ivl_27305 <= z2(17);
  tmp_ivl_27306 <= new_AGEMA_signal_3270 & tmp_ivl_27305;
  LPM_q_ivl_27309 <= tmp_ivl_27311 & tmp_ivl_27306;
  new_AGEMA_signal_3477 <= tmp_ivl_27313(1);
  n4193 <= tmp_ivl_27313(0);
  tmp_ivl_27313 <= LPM_d0_ivl_27317(0 + 1 downto 0);
  tmp_ivl_27319 <= z3(17);
  tmp_ivl_27320 <= new_AGEMA_signal_3527 & tmp_ivl_27319;
  LPM_q_ivl_27323 <= tmp_ivl_27325 & tmp_ivl_27320;
  tmp_ivl_27328 <= state_in_s1(233);
  tmp_ivl_27330 <= state_in_s0(233);
  tmp_ivl_27331 <= tmp_ivl_27328 & tmp_ivl_27330;
  LPM_q_ivl_27334 <= tmp_ivl_27336 & tmp_ivl_27331;
  new_AGEMA_signal_3788 <= tmp_ivl_27338(1);
  n3963 <= tmp_ivl_27338(0);
  tmp_ivl_27338 <= LPM_d0_ivl_27342(0 + 1 downto 0);
  tmp_ivl_27343 <= new_AGEMA_signal_3477 & n4193;
  LPM_q_ivl_27346 <= tmp_ivl_27348 & tmp_ivl_27343;
  tmp_ivl_27350 <= new_AGEMA_signal_3788 & n3963;
  LPM_q_ivl_27353 <= tmp_ivl_27355 & tmp_ivl_27350;
  new_AGEMA_signal_4102 <= tmp_ivl_27357(1);
  n4095 <= tmp_ivl_27357(0);
  tmp_ivl_27357 <= LPM_d0_ivl_27361(0 + 1 downto 0);
  tmp_ivl_27362 <= new_AGEMA_signal_4102 & n4095;
  LPM_q_ivl_27365 <= tmp_ivl_27367 & tmp_ivl_27362;
  tmp_ivl_27369 <= new_AGEMA_signal_4084 & n3987;
  LPM_q_ivl_27372 <= tmp_ivl_27374 & tmp_ivl_27369;
  new_AGEMA_signal_4391 <= tmp_ivl_27376(1);
  n3965 <= tmp_ivl_27376(0);
  tmp_ivl_27376 <= LPM_d0_ivl_27380(0 + 1 downto 0);
  tmp_ivl_27381 <= new_AGEMA_signal_2758 & n3265;
  LPM_q_ivl_27384 <= tmp_ivl_27386 & tmp_ivl_27381;
  tmp_ivl_27389 <= z2(34);
  tmp_ivl_27390 <= new_AGEMA_signal_3186 & tmp_ivl_27389;
  LPM_q_ivl_27393 <= tmp_ivl_27395 & tmp_ivl_27390;
  new_AGEMA_signal_3478 <= tmp_ivl_27397(1);
  n4159 <= tmp_ivl_27397(0);
  tmp_ivl_27397 <= LPM_d0_ivl_27401(0 + 1 downto 0);
  tmp_ivl_27403 <= z3(34);
  tmp_ivl_27404 <= new_AGEMA_signal_3546 & tmp_ivl_27403;
  LPM_q_ivl_27407 <= tmp_ivl_27409 & tmp_ivl_27404;
  tmp_ivl_27412 <= state_in_s1(218);
  tmp_ivl_27414 <= state_in_s0(218);
  tmp_ivl_27415 <= tmp_ivl_27412 & tmp_ivl_27414;
  LPM_q_ivl_27418 <= tmp_ivl_27420 & tmp_ivl_27415;
  new_AGEMA_signal_3789 <= tmp_ivl_27422(1);
  n3964 <= tmp_ivl_27422(0);
  tmp_ivl_27422 <= LPM_d0_ivl_27426(0 + 1 downto 0);
  tmp_ivl_27427 <= new_AGEMA_signal_3478 & n4159;
  LPM_q_ivl_27430 <= tmp_ivl_27432 & tmp_ivl_27427;
  tmp_ivl_27434 <= new_AGEMA_signal_3789 & n3964;
  LPM_q_ivl_27437 <= tmp_ivl_27439 & tmp_ivl_27434;
  new_AGEMA_signal_4103 <= tmp_ivl_27441(1);
  n4007 <= tmp_ivl_27441(0);
  tmp_ivl_27441 <= LPM_d0_ivl_27445(0 + 1 downto 0);
  tmp_ivl_27446 <= new_AGEMA_signal_4391 & n3965;
  LPM_q_ivl_27449 <= tmp_ivl_27451 & tmp_ivl_27446;
  tmp_ivl_27453 <= new_AGEMA_signal_4103 & n4007;
  LPM_q_ivl_27456 <= tmp_ivl_27458 & tmp_ivl_27453;
  tmp_ivl_27460 <= tmp_ivl_27464(1);
  tmp_ivl_27462 <= tmp_ivl_27464(0);
  tmp_ivl_27464 <= LPM_d0_ivl_27468(0 + 1 downto 0);
  tmp_ivl_27469 <= new_AGEMA_signal_2760 & n3281;
  LPM_q_ivl_27472 <= tmp_ivl_27474 & tmp_ivl_27469;
  tmp_ivl_27477 <= z2(18);
  tmp_ivl_27478 <= new_AGEMA_signal_3284 & tmp_ivl_27477;
  LPM_q_ivl_27481 <= tmp_ivl_27483 & tmp_ivl_27478;
  new_AGEMA_signal_3479 <= tmp_ivl_27485(1);
  n4191 <= tmp_ivl_27485(0);
  tmp_ivl_27485 <= LPM_d0_ivl_27489(0 + 1 downto 0);
  tmp_ivl_27491 <= z3(18);
  tmp_ivl_27492 <= new_AGEMA_signal_3528 & tmp_ivl_27491;
  LPM_q_ivl_27495 <= tmp_ivl_27497 & tmp_ivl_27492;
  tmp_ivl_27500 <= state_in_s1(234);
  tmp_ivl_27502 <= state_in_s0(234);
  tmp_ivl_27503 <= tmp_ivl_27500 & tmp_ivl_27502;
  LPM_q_ivl_27506 <= tmp_ivl_27508 & tmp_ivl_27503;
  new_AGEMA_signal_3790 <= tmp_ivl_27510(1);
  n3966 <= tmp_ivl_27510(0);
  tmp_ivl_27510 <= LPM_d0_ivl_27514(0 + 1 downto 0);
  tmp_ivl_27515 <= new_AGEMA_signal_3479 & n4191;
  LPM_q_ivl_27518 <= tmp_ivl_27520 & tmp_ivl_27515;
  tmp_ivl_27522 <= new_AGEMA_signal_3790 & n3966;
  LPM_q_ivl_27525 <= tmp_ivl_27527 & tmp_ivl_27522;
  new_AGEMA_signal_4104 <= tmp_ivl_27529(1);
  n4063 <= tmp_ivl_27529(0);
  tmp_ivl_27529 <= LPM_d0_ivl_27533(0 + 1 downto 0);
  tmp_ivl_27534 <= new_AGEMA_signal_2763 & n3264;
  LPM_q_ivl_27537 <= tmp_ivl_27539 & tmp_ivl_27534;
  tmp_ivl_27542 <= z2(35);
  tmp_ivl_27543 <= new_AGEMA_signal_3185 & tmp_ivl_27542;
  LPM_q_ivl_27546 <= tmp_ivl_27548 & tmp_ivl_27543;
  new_AGEMA_signal_3480 <= tmp_ivl_27550(1);
  n4157 <= tmp_ivl_27550(0);
  tmp_ivl_27550 <= LPM_d0_ivl_27554(0 + 1 downto 0);
  tmp_ivl_27556 <= z3(35);
  tmp_ivl_27557 <= new_AGEMA_signal_3547 & tmp_ivl_27556;
  LPM_q_ivl_27560 <= tmp_ivl_27562 & tmp_ivl_27557;
  tmp_ivl_27565 <= state_in_s1(219);
  tmp_ivl_27567 <= state_in_s0(219);
  tmp_ivl_27568 <= tmp_ivl_27565 & tmp_ivl_27567;
  LPM_q_ivl_27571 <= tmp_ivl_27573 & tmp_ivl_27568;
  new_AGEMA_signal_3791 <= tmp_ivl_27575(1);
  n3967 <= tmp_ivl_27575(0);
  tmp_ivl_27575 <= LPM_d0_ivl_27579(0 + 1 downto 0);
  tmp_ivl_27580 <= new_AGEMA_signal_3480 & n4157;
  LPM_q_ivl_27583 <= tmp_ivl_27585 & tmp_ivl_27580;
  tmp_ivl_27587 <= new_AGEMA_signal_3791 & n3967;
  LPM_q_ivl_27590 <= tmp_ivl_27592 & tmp_ivl_27587;
  new_AGEMA_signal_4105 <= tmp_ivl_27594(1);
  n4010 <= tmp_ivl_27594(0);
  tmp_ivl_27594 <= LPM_d0_ivl_27598(0 + 1 downto 0);
  tmp_ivl_27599 <= new_AGEMA_signal_4104 & n4063;
  LPM_q_ivl_27602 <= tmp_ivl_27604 & tmp_ivl_27599;
  tmp_ivl_27606 <= new_AGEMA_signal_4105 & n4010;
  LPM_q_ivl_27609 <= tmp_ivl_27611 & tmp_ivl_27606;
  new_AGEMA_signal_4392 <= tmp_ivl_27613(1);
  n3968 <= tmp_ivl_27613(0);
  tmp_ivl_27613 <= LPM_d0_ivl_27617(0 + 1 downto 0);
  tmp_ivl_27618 <= new_AGEMA_signal_4087 & n3989;
  LPM_q_ivl_27621 <= tmp_ivl_27623 & tmp_ivl_27618;
  tmp_ivl_27625 <= new_AGEMA_signal_4392 & n3968;
  LPM_q_ivl_27628 <= tmp_ivl_27630 & tmp_ivl_27625;
  tmp_ivl_27632 <= tmp_ivl_27636(1);
  tmp_ivl_27634 <= tmp_ivl_27636(0);
  tmp_ivl_27636 <= LPM_d0_ivl_27640(0 + 1 downto 0);
  tmp_ivl_27641 <= new_AGEMA_signal_4090 & n3992;
  LPM_q_ivl_27644 <= tmp_ivl_27646 & tmp_ivl_27641;
  tmp_ivl_27648 <= new_AGEMA_signal_4080 & n4076;
  LPM_q_ivl_27651 <= tmp_ivl_27653 & tmp_ivl_27648;
  new_AGEMA_signal_4393 <= tmp_ivl_27655(1);
  n3970 <= tmp_ivl_27655(0);
  tmp_ivl_27655 <= LPM_d0_ivl_27659(0 + 1 downto 0);
  tmp_ivl_27660 <= new_AGEMA_signal_2766 & n3263;
  LPM_q_ivl_27663 <= tmp_ivl_27665 & tmp_ivl_27660;
  tmp_ivl_27668 <= z2(36);
  tmp_ivl_27669 <= new_AGEMA_signal_3183 & tmp_ivl_27668;
  LPM_q_ivl_27672 <= tmp_ivl_27674 & tmp_ivl_27669;
  new_AGEMA_signal_3481 <= tmp_ivl_27676(1);
  n4155 <= tmp_ivl_27676(0);
  tmp_ivl_27676 <= LPM_d0_ivl_27680(0 + 1 downto 0);
  tmp_ivl_27682 <= z3(36);
  tmp_ivl_27683 <= new_AGEMA_signal_3548 & tmp_ivl_27682;
  LPM_q_ivl_27686 <= tmp_ivl_27688 & tmp_ivl_27683;
  tmp_ivl_27691 <= state_in_s1(220);
  tmp_ivl_27693 <= state_in_s0(220);
  tmp_ivl_27694 <= tmp_ivl_27691 & tmp_ivl_27693;
  LPM_q_ivl_27697 <= tmp_ivl_27699 & tmp_ivl_27694;
  new_AGEMA_signal_3792 <= tmp_ivl_27701(1);
  n3969 <= tmp_ivl_27701(0);
  tmp_ivl_27701 <= LPM_d0_ivl_27705(0 + 1 downto 0);
  tmp_ivl_27706 <= new_AGEMA_signal_3481 & n4155;
  LPM_q_ivl_27709 <= tmp_ivl_27711 & tmp_ivl_27706;
  tmp_ivl_27713 <= new_AGEMA_signal_3792 & n3969;
  LPM_q_ivl_27716 <= tmp_ivl_27718 & tmp_ivl_27713;
  new_AGEMA_signal_4106 <= tmp_ivl_27720(1);
  n4015 <= tmp_ivl_27720(0);
  tmp_ivl_27720 <= LPM_d0_ivl_27724(0 + 1 downto 0);
  tmp_ivl_27725 <= new_AGEMA_signal_4393 & n3970;
  LPM_q_ivl_27728 <= tmp_ivl_27730 & tmp_ivl_27725;
  tmp_ivl_27732 <= new_AGEMA_signal_4106 & n4015;
  LPM_q_ivl_27735 <= tmp_ivl_27737 & tmp_ivl_27732;
  tmp_ivl_27739 <= tmp_ivl_27743(1);
  tmp_ivl_27741 <= tmp_ivl_27743(0);
  tmp_ivl_27743 <= LPM_d0_ivl_27747(0 + 1 downto 0);
  tmp_ivl_27748 <= new_AGEMA_signal_4082 & n4264;
  LPM_q_ivl_27751 <= tmp_ivl_27753 & tmp_ivl_27748;
  tmp_ivl_27755 <= new_AGEMA_signal_4093 & n3996;
  LPM_q_ivl_27758 <= tmp_ivl_27760 & tmp_ivl_27755;
  new_AGEMA_signal_4394 <= tmp_ivl_27762(1);
  n3972 <= tmp_ivl_27762(0);
  tmp_ivl_27762 <= LPM_d0_ivl_27766(0 + 1 downto 0);
  tmp_ivl_27767 <= new_AGEMA_signal_2769 & n3262;
  LPM_q_ivl_27770 <= tmp_ivl_27772 & tmp_ivl_27767;
  tmp_ivl_27775 <= z2(37);
  tmp_ivl_27776 <= new_AGEMA_signal_3181 & tmp_ivl_27775;
  LPM_q_ivl_27779 <= tmp_ivl_27781 & tmp_ivl_27776;
  new_AGEMA_signal_3482 <= tmp_ivl_27783(1);
  n4153 <= tmp_ivl_27783(0);
  tmp_ivl_27783 <= LPM_d0_ivl_27787(0 + 1 downto 0);
  tmp_ivl_27789 <= z3(37);
  tmp_ivl_27790 <= new_AGEMA_signal_3549 & tmp_ivl_27789;
  LPM_q_ivl_27793 <= tmp_ivl_27795 & tmp_ivl_27790;
  tmp_ivl_27798 <= state_in_s1(221);
  tmp_ivl_27800 <= state_in_s0(221);
  tmp_ivl_27801 <= tmp_ivl_27798 & tmp_ivl_27800;
  LPM_q_ivl_27804 <= tmp_ivl_27806 & tmp_ivl_27801;
  new_AGEMA_signal_3793 <= tmp_ivl_27808(1);
  n3971 <= tmp_ivl_27808(0);
  tmp_ivl_27808 <= LPM_d0_ivl_27812(0 + 1 downto 0);
  tmp_ivl_27813 <= new_AGEMA_signal_3482 & n4153;
  LPM_q_ivl_27816 <= tmp_ivl_27818 & tmp_ivl_27813;
  tmp_ivl_27820 <= new_AGEMA_signal_3793 & n3971;
  LPM_q_ivl_27823 <= tmp_ivl_27825 & tmp_ivl_27820;
  new_AGEMA_signal_4107 <= tmp_ivl_27827(1);
  n4018 <= tmp_ivl_27827(0);
  tmp_ivl_27827 <= LPM_d0_ivl_27831(0 + 1 downto 0);
  tmp_ivl_27832 <= new_AGEMA_signal_4394 & n3972;
  LPM_q_ivl_27835 <= tmp_ivl_27837 & tmp_ivl_27832;
  tmp_ivl_27839 <= new_AGEMA_signal_4107 & n4018;
  LPM_q_ivl_27842 <= tmp_ivl_27844 & tmp_ivl_27839;
  tmp_ivl_27846 <= tmp_ivl_27850(1);
  tmp_ivl_27848 <= tmp_ivl_27850(0);
  tmp_ivl_27850 <= LPM_d0_ivl_27854(0 + 1 downto 0);
  tmp_ivl_27855 <= new_AGEMA_signal_4086 & n4254;
  LPM_q_ivl_27858 <= tmp_ivl_27860 & tmp_ivl_27855;
  tmp_ivl_27862 <= new_AGEMA_signal_4096 & n3998;
  LPM_q_ivl_27865 <= tmp_ivl_27867 & tmp_ivl_27862;
  new_AGEMA_signal_4395 <= tmp_ivl_27869(1);
  n3974 <= tmp_ivl_27869(0);
  tmp_ivl_27869 <= LPM_d0_ivl_27873(0 + 1 downto 0);
  tmp_ivl_27874 <= new_AGEMA_signal_2772 & n3261;
  LPM_q_ivl_27877 <= tmp_ivl_27879 & tmp_ivl_27874;
  tmp_ivl_27882 <= z2(38);
  tmp_ivl_27883 <= new_AGEMA_signal_3179 & tmp_ivl_27882;
  LPM_q_ivl_27886 <= tmp_ivl_27888 & tmp_ivl_27883;
  new_AGEMA_signal_3483 <= tmp_ivl_27890(1);
  n4151 <= tmp_ivl_27890(0);
  tmp_ivl_27890 <= LPM_d0_ivl_27894(0 + 1 downto 0);
  tmp_ivl_27896 <= z3(38);
  tmp_ivl_27897 <= new_AGEMA_signal_3550 & tmp_ivl_27896;
  LPM_q_ivl_27900 <= tmp_ivl_27902 & tmp_ivl_27897;
  tmp_ivl_27905 <= state_in_s1(222);
  tmp_ivl_27907 <= state_in_s0(222);
  tmp_ivl_27908 <= tmp_ivl_27905 & tmp_ivl_27907;
  LPM_q_ivl_27911 <= tmp_ivl_27913 & tmp_ivl_27908;
  new_AGEMA_signal_3794 <= tmp_ivl_27915(1);
  n3973 <= tmp_ivl_27915(0);
  tmp_ivl_27915 <= LPM_d0_ivl_27919(0 + 1 downto 0);
  tmp_ivl_27920 <= new_AGEMA_signal_3483 & n4151;
  LPM_q_ivl_27923 <= tmp_ivl_27925 & tmp_ivl_27920;
  tmp_ivl_27927 <= new_AGEMA_signal_3794 & n3973;
  LPM_q_ivl_27930 <= tmp_ivl_27932 & tmp_ivl_27927;
  new_AGEMA_signal_4108 <= tmp_ivl_27934(1);
  n4019 <= tmp_ivl_27934(0);
  tmp_ivl_27934 <= LPM_d0_ivl_27938(0 + 1 downto 0);
  tmp_ivl_27939 <= new_AGEMA_signal_4395 & n3974;
  LPM_q_ivl_27942 <= tmp_ivl_27944 & tmp_ivl_27939;
  tmp_ivl_27946 <= new_AGEMA_signal_4108 & n4019;
  LPM_q_ivl_27949 <= tmp_ivl_27951 & tmp_ivl_27946;
  tmp_ivl_27953 <= tmp_ivl_27957(1);
  tmp_ivl_27955 <= tmp_ivl_27957(0);
  tmp_ivl_27957 <= LPM_d0_ivl_27961(0 + 1 downto 0);
  tmp_ivl_27962 <= new_AGEMA_signal_4089 & n4241;
  LPM_q_ivl_27965 <= tmp_ivl_27967 & tmp_ivl_27962;
  tmp_ivl_27969 <= new_AGEMA_signal_4099 & n4002;
  LPM_q_ivl_27972 <= tmp_ivl_27974 & tmp_ivl_27969;
  new_AGEMA_signal_4396 <= tmp_ivl_27976(1);
  n3976 <= tmp_ivl_27976(0);
  tmp_ivl_27976 <= LPM_d0_ivl_27980(0 + 1 downto 0);
  tmp_ivl_27981 <= new_AGEMA_signal_2775 & n3260;
  LPM_q_ivl_27984 <= tmp_ivl_27986 & tmp_ivl_27981;
  tmp_ivl_27989 <= z2(39);
  tmp_ivl_27990 <= new_AGEMA_signal_3176 & tmp_ivl_27989;
  LPM_q_ivl_27993 <= tmp_ivl_27995 & tmp_ivl_27990;
  new_AGEMA_signal_3484 <= tmp_ivl_27997(1);
  n4149 <= tmp_ivl_27997(0);
  tmp_ivl_27997 <= LPM_d0_ivl_28001(0 + 1 downto 0);
  tmp_ivl_28003 <= z3(39);
  tmp_ivl_28004 <= new_AGEMA_signal_3551 & tmp_ivl_28003;
  LPM_q_ivl_28007 <= tmp_ivl_28009 & tmp_ivl_28004;
  tmp_ivl_28012 <= state_in_s1(223);
  tmp_ivl_28014 <= state_in_s0(223);
  tmp_ivl_28015 <= tmp_ivl_28012 & tmp_ivl_28014;
  LPM_q_ivl_28018 <= tmp_ivl_28020 & tmp_ivl_28015;
  new_AGEMA_signal_3795 <= tmp_ivl_28022(1);
  n3975 <= tmp_ivl_28022(0);
  tmp_ivl_28022 <= LPM_d0_ivl_28026(0 + 1 downto 0);
  tmp_ivl_28027 <= new_AGEMA_signal_3484 & n4149;
  LPM_q_ivl_28030 <= tmp_ivl_28032 & tmp_ivl_28027;
  tmp_ivl_28034 <= new_AGEMA_signal_3795 & n3975;
  LPM_q_ivl_28037 <= tmp_ivl_28039 & tmp_ivl_28034;
  new_AGEMA_signal_4109 <= tmp_ivl_28041(1);
  n4023 <= tmp_ivl_28041(0);
  tmp_ivl_28041 <= LPM_d0_ivl_28045(0 + 1 downto 0);
  tmp_ivl_28046 <= new_AGEMA_signal_4396 & n3976;
  LPM_q_ivl_28049 <= tmp_ivl_28051 & tmp_ivl_28046;
  tmp_ivl_28053 <= new_AGEMA_signal_4109 & n4023;
  LPM_q_ivl_28056 <= tmp_ivl_28058 & tmp_ivl_28053;
  tmp_ivl_28060 <= tmp_ivl_28064(1);
  tmp_ivl_28062 <= tmp_ivl_28064(0);
  tmp_ivl_28064 <= LPM_d0_ivl_28068(0 + 1 downto 0);
  tmp_ivl_28069 <= new_AGEMA_signal_4091 & n4230;
  LPM_q_ivl_28072 <= tmp_ivl_28074 & tmp_ivl_28069;
  tmp_ivl_28076 <= new_AGEMA_signal_4101 & n4006;
  LPM_q_ivl_28079 <= tmp_ivl_28081 & tmp_ivl_28076;
  new_AGEMA_signal_4397 <= tmp_ivl_28083(1);
  n3978 <= tmp_ivl_28083(0);
  tmp_ivl_28083 <= LPM_d0_ivl_28087(0 + 1 downto 0);
  tmp_ivl_28088 <= new_AGEMA_signal_2778 & n3259;
  LPM_q_ivl_28091 <= tmp_ivl_28093 & tmp_ivl_28088;
  tmp_ivl_28096 <= z2(40);
  tmp_ivl_28097 <= new_AGEMA_signal_3177 & tmp_ivl_28096;
  LPM_q_ivl_28100 <= tmp_ivl_28102 & tmp_ivl_28097;
  new_AGEMA_signal_3485 <= tmp_ivl_28104(1);
  n4147 <= tmp_ivl_28104(0);
  tmp_ivl_28104 <= LPM_d0_ivl_28108(0 + 1 downto 0);
  tmp_ivl_28110 <= z3(40);
  tmp_ivl_28111 <= new_AGEMA_signal_3553 & tmp_ivl_28110;
  LPM_q_ivl_28114 <= tmp_ivl_28116 & tmp_ivl_28111;
  tmp_ivl_28119 <= state_in_s1(208);
  tmp_ivl_28121 <= state_in_s0(208);
  tmp_ivl_28122 <= tmp_ivl_28119 & tmp_ivl_28121;
  LPM_q_ivl_28125 <= tmp_ivl_28127 & tmp_ivl_28122;
  new_AGEMA_signal_3796 <= tmp_ivl_28129(1);
  n3977 <= tmp_ivl_28129(0);
  tmp_ivl_28129 <= LPM_d0_ivl_28133(0 + 1 downto 0);
  tmp_ivl_28134 <= new_AGEMA_signal_3485 & n4147;
  LPM_q_ivl_28137 <= tmp_ivl_28139 & tmp_ivl_28134;
  tmp_ivl_28141 <= new_AGEMA_signal_3796 & n3977;
  LPM_q_ivl_28144 <= tmp_ivl_28146 & tmp_ivl_28141;
  new_AGEMA_signal_4110 <= tmp_ivl_28148(1);
  n4027 <= tmp_ivl_28148(0);
  tmp_ivl_28148 <= LPM_d0_ivl_28152(0 + 1 downto 0);
  tmp_ivl_28153 <= new_AGEMA_signal_4397 & n3978;
  LPM_q_ivl_28156 <= tmp_ivl_28158 & tmp_ivl_28153;
  tmp_ivl_28160 <= new_AGEMA_signal_4110 & n4027;
  LPM_q_ivl_28163 <= tmp_ivl_28165 & tmp_ivl_28160;
  tmp_ivl_28167 <= tmp_ivl_28171(1);
  tmp_ivl_28169 <= tmp_ivl_28171(0);
  tmp_ivl_28171 <= LPM_d0_ivl_28175(0 + 1 downto 0);
  tmp_ivl_28176 <= new_AGEMA_signal_4095 & n4094;
  LPM_q_ivl_28179 <= tmp_ivl_28181 & tmp_ivl_28176;
  tmp_ivl_28183 <= new_AGEMA_signal_4103 & n4007;
  LPM_q_ivl_28186 <= tmp_ivl_28188 & tmp_ivl_28183;
  new_AGEMA_signal_4398 <= tmp_ivl_28190(1);
  n3980 <= tmp_ivl_28190(0);
  tmp_ivl_28190 <= LPM_d0_ivl_28194(0 + 1 downto 0);
  tmp_ivl_28195 <= new_AGEMA_signal_2780 & n3258;
  LPM_q_ivl_28198 <= tmp_ivl_28200 & tmp_ivl_28195;
  tmp_ivl_28203 <= z2(41);
  tmp_ivl_28204 <= new_AGEMA_signal_3184 & tmp_ivl_28203;
  LPM_q_ivl_28207 <= tmp_ivl_28209 & tmp_ivl_28204;
  new_AGEMA_signal_3486 <= tmp_ivl_28211(1);
  n4145 <= tmp_ivl_28211(0);
  tmp_ivl_28211 <= LPM_d0_ivl_28215(0 + 1 downto 0);
  tmp_ivl_28217 <= z3(41);
  tmp_ivl_28218 <= new_AGEMA_signal_3554 & tmp_ivl_28217;
  LPM_q_ivl_28221 <= tmp_ivl_28223 & tmp_ivl_28218;
  tmp_ivl_28226 <= state_in_s1(209);
  tmp_ivl_28228 <= state_in_s0(209);
  tmp_ivl_28229 <= tmp_ivl_28226 & tmp_ivl_28228;
  LPM_q_ivl_28232 <= tmp_ivl_28234 & tmp_ivl_28229;
  new_AGEMA_signal_3797 <= tmp_ivl_28236(1);
  n3979 <= tmp_ivl_28236(0);
  tmp_ivl_28236 <= LPM_d0_ivl_28240(0 + 1 downto 0);
  tmp_ivl_28241 <= new_AGEMA_signal_3486 & n4145;
  LPM_q_ivl_28244 <= tmp_ivl_28246 & tmp_ivl_28241;
  tmp_ivl_28248 <= new_AGEMA_signal_3797 & n3979;
  LPM_q_ivl_28251 <= tmp_ivl_28253 & tmp_ivl_28248;
  new_AGEMA_signal_4111 <= tmp_ivl_28255(1);
  n4029 <= tmp_ivl_28255(0);
  tmp_ivl_28255 <= LPM_d0_ivl_28259(0 + 1 downto 0);
  tmp_ivl_28260 <= new_AGEMA_signal_4398 & n3980;
  LPM_q_ivl_28263 <= tmp_ivl_28265 & tmp_ivl_28260;
  tmp_ivl_28267 <= new_AGEMA_signal_4111 & n4029;
  LPM_q_ivl_28270 <= tmp_ivl_28272 & tmp_ivl_28267;
  tmp_ivl_28274 <= tmp_ivl_28278(1);
  tmp_ivl_28276 <= tmp_ivl_28278(0);
  tmp_ivl_28278 <= LPM_d0_ivl_28282(0 + 1 downto 0);
  tmp_ivl_28283 <= new_AGEMA_signal_4098 & n4044;
  LPM_q_ivl_28286 <= tmp_ivl_28288 & tmp_ivl_28283;
  tmp_ivl_28290 <= new_AGEMA_signal_4105 & n4010;
  LPM_q_ivl_28293 <= tmp_ivl_28295 & tmp_ivl_28290;
  new_AGEMA_signal_4399 <= tmp_ivl_28297(1);
  n3982 <= tmp_ivl_28297(0);
  tmp_ivl_28297 <= LPM_d0_ivl_28301(0 + 1 downto 0);
  tmp_ivl_28302 <= new_AGEMA_signal_2783 & n3257;
  LPM_q_ivl_28305 <= tmp_ivl_28307 & tmp_ivl_28302;
  tmp_ivl_28310 <= z2(42);
  tmp_ivl_28311 <= new_AGEMA_signal_3182 & tmp_ivl_28310;
  LPM_q_ivl_28314 <= tmp_ivl_28316 & tmp_ivl_28311;
  new_AGEMA_signal_3487 <= tmp_ivl_28318(1);
  n4143 <= tmp_ivl_28318(0);
  tmp_ivl_28318 <= LPM_d0_ivl_28322(0 + 1 downto 0);
  tmp_ivl_28324 <= z3(42);
  tmp_ivl_28325 <= new_AGEMA_signal_3555 & tmp_ivl_28324;
  LPM_q_ivl_28328 <= tmp_ivl_28330 & tmp_ivl_28325;
  tmp_ivl_28333 <= state_in_s1(210);
  tmp_ivl_28335 <= state_in_s0(210);
  tmp_ivl_28336 <= tmp_ivl_28333 & tmp_ivl_28335;
  LPM_q_ivl_28339 <= tmp_ivl_28341 & tmp_ivl_28336;
  new_AGEMA_signal_3798 <= tmp_ivl_28343(1);
  n3981 <= tmp_ivl_28343(0);
  tmp_ivl_28343 <= LPM_d0_ivl_28347(0 + 1 downto 0);
  tmp_ivl_28348 <= new_AGEMA_signal_3487 & n4143;
  LPM_q_ivl_28351 <= tmp_ivl_28353 & tmp_ivl_28348;
  tmp_ivl_28355 <= new_AGEMA_signal_3798 & n3981;
  LPM_q_ivl_28358 <= tmp_ivl_28360 & tmp_ivl_28355;
  new_AGEMA_signal_4112 <= tmp_ivl_28362(1);
  n4032 <= tmp_ivl_28362(0);
  tmp_ivl_28362 <= LPM_d0_ivl_28366(0 + 1 downto 0);
  tmp_ivl_28367 <= new_AGEMA_signal_4399 & n3982;
  LPM_q_ivl_28370 <= tmp_ivl_28372 & tmp_ivl_28367;
  tmp_ivl_28374 <= new_AGEMA_signal_4112 & n4032;
  LPM_q_ivl_28377 <= tmp_ivl_28379 & tmp_ivl_28374;
  tmp_ivl_28381 <= tmp_ivl_28385(1);
  tmp_ivl_28383 <= tmp_ivl_28385(0);
  tmp_ivl_28385 <= LPM_d0_ivl_28389(0 + 1 downto 0);
  tmp_ivl_28390 <= new_AGEMA_signal_2786 & n3256;
  LPM_q_ivl_28393 <= tmp_ivl_28395 & tmp_ivl_28390;
  tmp_ivl_28398 <= z2(43);
  tmp_ivl_28399 <= new_AGEMA_signal_3180 & tmp_ivl_28398;
  LPM_q_ivl_28402 <= tmp_ivl_28404 & tmp_ivl_28399;
  new_AGEMA_signal_3488 <= tmp_ivl_28406(1);
  n4141 <= tmp_ivl_28406(0);
  tmp_ivl_28406 <= LPM_d0_ivl_28410(0 + 1 downto 0);
  tmp_ivl_28412 <= z3(43);
  tmp_ivl_28413 <= new_AGEMA_signal_3556 & tmp_ivl_28412;
  LPM_q_ivl_28416 <= tmp_ivl_28418 & tmp_ivl_28413;
  tmp_ivl_28421 <= state_in_s1(211);
  tmp_ivl_28423 <= state_in_s0(211);
  tmp_ivl_28424 <= tmp_ivl_28421 & tmp_ivl_28423;
  LPM_q_ivl_28427 <= tmp_ivl_28429 & tmp_ivl_28424;
  new_AGEMA_signal_3799 <= tmp_ivl_28431(1);
  n3983 <= tmp_ivl_28431(0);
  tmp_ivl_28431 <= LPM_d0_ivl_28435(0 + 1 downto 0);
  tmp_ivl_28436 <= new_AGEMA_signal_3488 & n4141;
  LPM_q_ivl_28439 <= tmp_ivl_28441 & tmp_ivl_28436;
  tmp_ivl_28443 <= new_AGEMA_signal_3799 & n3983;
  LPM_q_ivl_28446 <= tmp_ivl_28448 & tmp_ivl_28443;
  new_AGEMA_signal_4113 <= tmp_ivl_28450(1);
  n4035 <= tmp_ivl_28450(0);
  tmp_ivl_28450 <= LPM_d0_ivl_28454(0 + 1 downto 0);
  tmp_ivl_28455 <= new_AGEMA_signal_4113 & n4035;
  LPM_q_ivl_28458 <= tmp_ivl_28460 & tmp_ivl_28455;
  tmp_ivl_28462 <= new_AGEMA_signal_4081 & n3984;
  LPM_q_ivl_28465 <= tmp_ivl_28467 & tmp_ivl_28462;
  new_AGEMA_signal_4400 <= tmp_ivl_28469(1);
  n3985 <= tmp_ivl_28469(0);
  tmp_ivl_28469 <= LPM_d0_ivl_28473(0 + 1 downto 0);
  tmp_ivl_28474 <= new_AGEMA_signal_4400 & n3985;
  LPM_q_ivl_28477 <= tmp_ivl_28479 & tmp_ivl_28474;
  tmp_ivl_28481 <= new_AGEMA_signal_4106 & n4015;
  LPM_q_ivl_28484 <= tmp_ivl_28486 & tmp_ivl_28481;
  tmp_ivl_28488 <= tmp_ivl_28492(1);
  tmp_ivl_28490 <= tmp_ivl_28492(0);
  tmp_ivl_28492 <= LPM_d0_ivl_28496(0 + 1 downto 0);
  tmp_ivl_28497 <= new_AGEMA_signal_2788 & n3255;
  LPM_q_ivl_28500 <= tmp_ivl_28502 & tmp_ivl_28497;
  tmp_ivl_28505 <= z2(44);
  tmp_ivl_28506 <= new_AGEMA_signal_3178 & tmp_ivl_28505;
  LPM_q_ivl_28509 <= tmp_ivl_28511 & tmp_ivl_28506;
  new_AGEMA_signal_3489 <= tmp_ivl_28513(1);
  n4139 <= tmp_ivl_28513(0);
  tmp_ivl_28513 <= LPM_d0_ivl_28517(0 + 1 downto 0);
  tmp_ivl_28519 <= z3(44);
  tmp_ivl_28520 <= new_AGEMA_signal_3557 & tmp_ivl_28519;
  LPM_q_ivl_28523 <= tmp_ivl_28525 & tmp_ivl_28520;
  tmp_ivl_28528 <= state_in_s1(212);
  tmp_ivl_28530 <= state_in_s0(212);
  tmp_ivl_28531 <= tmp_ivl_28528 & tmp_ivl_28530;
  LPM_q_ivl_28534 <= tmp_ivl_28536 & tmp_ivl_28531;
  new_AGEMA_signal_3800 <= tmp_ivl_28538(1);
  n3986 <= tmp_ivl_28538(0);
  tmp_ivl_28538 <= LPM_d0_ivl_28542(0 + 1 downto 0);
  tmp_ivl_28543 <= new_AGEMA_signal_3489 & n4139;
  LPM_q_ivl_28546 <= tmp_ivl_28548 & tmp_ivl_28543;
  tmp_ivl_28550 <= new_AGEMA_signal_3800 & n3986;
  LPM_q_ivl_28553 <= tmp_ivl_28555 & tmp_ivl_28550;
  new_AGEMA_signal_4114 <= tmp_ivl_28557(1);
  n4046 <= tmp_ivl_28557(0);
  tmp_ivl_28557 <= LPM_d0_ivl_28561(0 + 1 downto 0);
  tmp_ivl_28562 <= new_AGEMA_signal_4114 & n4046;
  LPM_q_ivl_28565 <= tmp_ivl_28567 & tmp_ivl_28562;
  tmp_ivl_28569 <= new_AGEMA_signal_4084 & n3987;
  LPM_q_ivl_28572 <= tmp_ivl_28574 & tmp_ivl_28569;
  new_AGEMA_signal_4401 <= tmp_ivl_28576(1);
  n3988 <= tmp_ivl_28576(0);
  tmp_ivl_28576 <= LPM_d0_ivl_28580(0 + 1 downto 0);
  tmp_ivl_28581 <= new_AGEMA_signal_4401 & n3988;
  LPM_q_ivl_28584 <= tmp_ivl_28586 & tmp_ivl_28581;
  tmp_ivl_28588 <= new_AGEMA_signal_4107 & n4018;
  LPM_q_ivl_28591 <= tmp_ivl_28593 & tmp_ivl_28588;
  tmp_ivl_28595 <= tmp_ivl_28599(1);
  tmp_ivl_28597 <= tmp_ivl_28599(0);
  tmp_ivl_28599 <= LPM_d0_ivl_28603(0 + 1 downto 0);
  tmp_ivl_28604 <= new_AGEMA_signal_4087 & n3989;
  LPM_q_ivl_28607 <= tmp_ivl_28609 & tmp_ivl_28604;
  tmp_ivl_28611 <= new_AGEMA_signal_4108 & n4019;
  LPM_q_ivl_28614 <= tmp_ivl_28616 & tmp_ivl_28611;
  new_AGEMA_signal_4402 <= tmp_ivl_28618(1);
  n3991 <= tmp_ivl_28618(0);
  tmp_ivl_28618 <= LPM_d0_ivl_28622(0 + 1 downto 0);
  tmp_ivl_28623 <= new_AGEMA_signal_2790 & n3254;
  LPM_q_ivl_28626 <= tmp_ivl_28628 & tmp_ivl_28623;
  tmp_ivl_28631 <= z2(45);
  tmp_ivl_28632 <= new_AGEMA_signal_3175 & tmp_ivl_28631;
  LPM_q_ivl_28635 <= tmp_ivl_28637 & tmp_ivl_28632;
  new_AGEMA_signal_3490 <= tmp_ivl_28639(1);
  n4137 <= tmp_ivl_28639(0);
  tmp_ivl_28639 <= LPM_d0_ivl_28643(0 + 1 downto 0);
  tmp_ivl_28645 <= z3(45);
  tmp_ivl_28646 <= new_AGEMA_signal_3558 & tmp_ivl_28645;
  LPM_q_ivl_28649 <= tmp_ivl_28651 & tmp_ivl_28646;
  tmp_ivl_28654 <= state_in_s1(213);
  tmp_ivl_28656 <= state_in_s0(213);
  tmp_ivl_28657 <= tmp_ivl_28654 & tmp_ivl_28656;
  LPM_q_ivl_28660 <= tmp_ivl_28662 & tmp_ivl_28657;
  new_AGEMA_signal_3801 <= tmp_ivl_28664(1);
  n3990 <= tmp_ivl_28664(0);
  tmp_ivl_28664 <= LPM_d0_ivl_28668(0 + 1 downto 0);
  tmp_ivl_28669 <= new_AGEMA_signal_3490 & n4137;
  LPM_q_ivl_28672 <= tmp_ivl_28674 & tmp_ivl_28669;
  tmp_ivl_28676 <= new_AGEMA_signal_3801 & n3990;
  LPM_q_ivl_28679 <= tmp_ivl_28681 & tmp_ivl_28676;
  new_AGEMA_signal_4115 <= tmp_ivl_28683(1);
  n4050 <= tmp_ivl_28683(0);
  tmp_ivl_28683 <= LPM_d0_ivl_28687(0 + 1 downto 0);
  tmp_ivl_28688 <= new_AGEMA_signal_4402 & n3991;
  LPM_q_ivl_28691 <= tmp_ivl_28693 & tmp_ivl_28688;
  tmp_ivl_28695 <= new_AGEMA_signal_4115 & n4050;
  LPM_q_ivl_28698 <= tmp_ivl_28700 & tmp_ivl_28695;
  tmp_ivl_28702 <= tmp_ivl_28706(1);
  tmp_ivl_28704 <= tmp_ivl_28706(0);
  tmp_ivl_28706 <= LPM_d0_ivl_28710(0 + 1 downto 0);
  tmp_ivl_28711 <= new_AGEMA_signal_4090 & n3992;
  LPM_q_ivl_28714 <= tmp_ivl_28716 & tmp_ivl_28711;
  tmp_ivl_28718 <= new_AGEMA_signal_4109 & n4023;
  LPM_q_ivl_28721 <= tmp_ivl_28723 & tmp_ivl_28718;
  new_AGEMA_signal_4403 <= tmp_ivl_28725(1);
  n3994 <= tmp_ivl_28725(0);
  tmp_ivl_28725 <= LPM_d0_ivl_28729(0 + 1 downto 0);
  tmp_ivl_28730 <= new_AGEMA_signal_2793 & n3253;
  LPM_q_ivl_28733 <= tmp_ivl_28735 & tmp_ivl_28730;
  tmp_ivl_28738 <= z2(46);
  tmp_ivl_28739 <= new_AGEMA_signal_3193 & tmp_ivl_28738;
  LPM_q_ivl_28742 <= tmp_ivl_28744 & tmp_ivl_28739;
  new_AGEMA_signal_3491 <= tmp_ivl_28746(1);
  n4135 <= tmp_ivl_28746(0);
  tmp_ivl_28746 <= LPM_d0_ivl_28750(0 + 1 downto 0);
  tmp_ivl_28752 <= z3(46);
  tmp_ivl_28753 <= new_AGEMA_signal_3559 & tmp_ivl_28752;
  LPM_q_ivl_28756 <= tmp_ivl_28758 & tmp_ivl_28753;
  tmp_ivl_28761 <= state_in_s1(214);
  tmp_ivl_28763 <= state_in_s0(214);
  tmp_ivl_28764 <= tmp_ivl_28761 & tmp_ivl_28763;
  LPM_q_ivl_28767 <= tmp_ivl_28769 & tmp_ivl_28764;
  new_AGEMA_signal_3802 <= tmp_ivl_28771(1);
  n3993 <= tmp_ivl_28771(0);
  tmp_ivl_28771 <= LPM_d0_ivl_28775(0 + 1 downto 0);
  tmp_ivl_28776 <= new_AGEMA_signal_3491 & n4135;
  LPM_q_ivl_28779 <= tmp_ivl_28781 & tmp_ivl_28776;
  tmp_ivl_28783 <= new_AGEMA_signal_3802 & n3993;
  LPM_q_ivl_28786 <= tmp_ivl_28788 & tmp_ivl_28783;
  new_AGEMA_signal_4116 <= tmp_ivl_28790(1);
  n4055 <= tmp_ivl_28790(0);
  tmp_ivl_28790 <= LPM_d0_ivl_28794(0 + 1 downto 0);
  tmp_ivl_28795 <= new_AGEMA_signal_4403 & n3994;
  LPM_q_ivl_28798 <= tmp_ivl_28800 & tmp_ivl_28795;
  tmp_ivl_28802 <= new_AGEMA_signal_4116 & n4055;
  LPM_q_ivl_28805 <= tmp_ivl_28807 & tmp_ivl_28802;
  tmp_ivl_28809 <= tmp_ivl_28813(1);
  tmp_ivl_28811 <= tmp_ivl_28813(0);
  tmp_ivl_28813 <= LPM_d0_ivl_28817(0 + 1 downto 0);
  tmp_ivl_28818 <= new_AGEMA_signal_2795 & n3252;
  LPM_q_ivl_28821 <= tmp_ivl_28823 & tmp_ivl_28818;
  tmp_ivl_28826 <= z2(47);
  tmp_ivl_28827 <= new_AGEMA_signal_3191 & tmp_ivl_28826;
  LPM_q_ivl_28830 <= tmp_ivl_28832 & tmp_ivl_28827;
  new_AGEMA_signal_3492 <= tmp_ivl_28834(1);
  n4133 <= tmp_ivl_28834(0);
  tmp_ivl_28834 <= LPM_d0_ivl_28838(0 + 1 downto 0);
  tmp_ivl_28840 <= z3(47);
  tmp_ivl_28841 <= new_AGEMA_signal_3560 & tmp_ivl_28840;
  LPM_q_ivl_28844 <= tmp_ivl_28846 & tmp_ivl_28841;
  tmp_ivl_28849 <= state_in_s1(215);
  tmp_ivl_28851 <= state_in_s0(215);
  tmp_ivl_28852 <= tmp_ivl_28849 & tmp_ivl_28851;
  LPM_q_ivl_28855 <= tmp_ivl_28857 & tmp_ivl_28852;
  new_AGEMA_signal_3803 <= tmp_ivl_28859(1);
  n3995 <= tmp_ivl_28859(0);
  tmp_ivl_28859 <= LPM_d0_ivl_28863(0 + 1 downto 0);
  tmp_ivl_28864 <= new_AGEMA_signal_3492 & n4133;
  LPM_q_ivl_28867 <= tmp_ivl_28869 & tmp_ivl_28864;
  tmp_ivl_28871 <= new_AGEMA_signal_3803 & n3995;
  LPM_q_ivl_28874 <= tmp_ivl_28876 & tmp_ivl_28871;
  new_AGEMA_signal_4117 <= tmp_ivl_28878(1);
  n4038 <= tmp_ivl_28878(0);
  tmp_ivl_28878 <= LPM_d0_ivl_28882(0 + 1 downto 0);
  tmp_ivl_28883 <= new_AGEMA_signal_4117 & n4038;
  LPM_q_ivl_28886 <= tmp_ivl_28888 & tmp_ivl_28883;
  tmp_ivl_28890 <= new_AGEMA_signal_4093 & n3996;
  LPM_q_ivl_28893 <= tmp_ivl_28895 & tmp_ivl_28890;
  new_AGEMA_signal_4404 <= tmp_ivl_28897(1);
  n3997 <= tmp_ivl_28897(0);
  tmp_ivl_28897 <= LPM_d0_ivl_28901(0 + 1 downto 0);
  tmp_ivl_28902 <= new_AGEMA_signal_4404 & n3997;
  LPM_q_ivl_28905 <= tmp_ivl_28907 & tmp_ivl_28902;
  tmp_ivl_28909 <= new_AGEMA_signal_4110 & n4027;
  LPM_q_ivl_28912 <= tmp_ivl_28914 & tmp_ivl_28909;
  tmp_ivl_28916 <= tmp_ivl_28920(1);
  tmp_ivl_28918 <= tmp_ivl_28920(0);
  tmp_ivl_28920 <= LPM_d0_ivl_28924(0 + 1 downto 0);
  tmp_ivl_28925 <= new_AGEMA_signal_4096 & n3998;
  LPM_q_ivl_28928 <= tmp_ivl_28930 & tmp_ivl_28925;
  tmp_ivl_28932 <= new_AGEMA_signal_4111 & n4029;
  LPM_q_ivl_28935 <= tmp_ivl_28937 & tmp_ivl_28932;
  new_AGEMA_signal_4405 <= tmp_ivl_28939(1);
  n4000 <= tmp_ivl_28939(0);
  tmp_ivl_28939 <= LPM_d0_ivl_28943(0 + 1 downto 0);
  tmp_ivl_28944 <= new_AGEMA_signal_2797 & n3251;
  LPM_q_ivl_28947 <= tmp_ivl_28949 & tmp_ivl_28944;
  tmp_ivl_28952 <= z2(48);
  tmp_ivl_28953 <= new_AGEMA_signal_3189 & tmp_ivl_28952;
  LPM_q_ivl_28956 <= tmp_ivl_28958 & tmp_ivl_28953;
  new_AGEMA_signal_3493 <= tmp_ivl_28960(1);
  n4131 <= tmp_ivl_28960(0);
  tmp_ivl_28960 <= LPM_d0_ivl_28964(0 + 1 downto 0);
  tmp_ivl_28966 <= z3(48);
  tmp_ivl_28967 <= new_AGEMA_signal_3561 & tmp_ivl_28966;
  LPM_q_ivl_28970 <= tmp_ivl_28972 & tmp_ivl_28967;
  tmp_ivl_28975 <= state_in_s1(200);
  tmp_ivl_28977 <= state_in_s0(200);
  tmp_ivl_28978 <= tmp_ivl_28975 & tmp_ivl_28977;
  LPM_q_ivl_28981 <= tmp_ivl_28983 & tmp_ivl_28978;
  new_AGEMA_signal_3804 <= tmp_ivl_28985(1);
  n3999 <= tmp_ivl_28985(0);
  tmp_ivl_28985 <= LPM_d0_ivl_28989(0 + 1 downto 0);
  tmp_ivl_28990 <= new_AGEMA_signal_3493 & n4131;
  LPM_q_ivl_28993 <= tmp_ivl_28995 & tmp_ivl_28990;
  tmp_ivl_28997 <= new_AGEMA_signal_3804 & n3999;
  LPM_q_ivl_29000 <= tmp_ivl_29002 & tmp_ivl_28997;
  new_AGEMA_signal_4118 <= tmp_ivl_29004(1);
  n4058 <= tmp_ivl_29004(0);
  tmp_ivl_29004 <= LPM_d0_ivl_29008(0 + 1 downto 0);
  tmp_ivl_29009 <= new_AGEMA_signal_4405 & n4000;
  LPM_q_ivl_29012 <= tmp_ivl_29014 & tmp_ivl_29009;
  tmp_ivl_29016 <= new_AGEMA_signal_4118 & n4058;
  LPM_q_ivl_29019 <= tmp_ivl_29021 & tmp_ivl_29016;
  tmp_ivl_29023 <= tmp_ivl_29027(1);
  tmp_ivl_29025 <= tmp_ivl_29027(0);
  tmp_ivl_29027 <= LPM_d0_ivl_29031(0 + 1 downto 0);
  tmp_ivl_29032 <= new_AGEMA_signal_2800 & n3250;
  LPM_q_ivl_29035 <= tmp_ivl_29037 & tmp_ivl_29032;
  tmp_ivl_29040 <= z2(49);
  tmp_ivl_29041 <= new_AGEMA_signal_3196 & tmp_ivl_29040;
  LPM_q_ivl_29044 <= tmp_ivl_29046 & tmp_ivl_29041;
  new_AGEMA_signal_3494 <= tmp_ivl_29048(1);
  n4128 <= tmp_ivl_29048(0);
  tmp_ivl_29048 <= LPM_d0_ivl_29052(0 + 1 downto 0);
  tmp_ivl_29054 <= z3(49);
  tmp_ivl_29055 <= new_AGEMA_signal_3562 & tmp_ivl_29054;
  LPM_q_ivl_29058 <= tmp_ivl_29060 & tmp_ivl_29055;
  tmp_ivl_29063 <= state_in_s1(201);
  tmp_ivl_29065 <= state_in_s0(201);
  tmp_ivl_29066 <= tmp_ivl_29063 & tmp_ivl_29065;
  LPM_q_ivl_29069 <= tmp_ivl_29071 & tmp_ivl_29066;
  new_AGEMA_signal_3805 <= tmp_ivl_29073(1);
  n4001 <= tmp_ivl_29073(0);
  tmp_ivl_29073 <= LPM_d0_ivl_29077(0 + 1 downto 0);
  tmp_ivl_29078 <= new_AGEMA_signal_3494 & n4128;
  LPM_q_ivl_29081 <= tmp_ivl_29083 & tmp_ivl_29078;
  tmp_ivl_29085 <= new_AGEMA_signal_3805 & n4001;
  LPM_q_ivl_29088 <= tmp_ivl_29090 & tmp_ivl_29085;
  new_AGEMA_signal_4119 <= tmp_ivl_29092(1);
  n4074 <= tmp_ivl_29092(0);
  tmp_ivl_29092 <= LPM_d0_ivl_29096(0 + 1 downto 0);
  tmp_ivl_29097 <= new_AGEMA_signal_4099 & n4002;
  LPM_q_ivl_29100 <= tmp_ivl_29102 & tmp_ivl_29097;
  tmp_ivl_29104 <= new_AGEMA_signal_4112 & n4032;
  LPM_q_ivl_29107 <= tmp_ivl_29109 & tmp_ivl_29104;
  new_AGEMA_signal_4406 <= tmp_ivl_29111(1);
  n4003 <= tmp_ivl_29111(0);
  tmp_ivl_29111 <= LPM_d0_ivl_29115(0 + 1 downto 0);
  tmp_ivl_29116 <= new_AGEMA_signal_4119 & n4074;
  LPM_q_ivl_29119 <= tmp_ivl_29121 & tmp_ivl_29116;
  tmp_ivl_29123 <= new_AGEMA_signal_4406 & n4003;
  LPM_q_ivl_29126 <= tmp_ivl_29128 & tmp_ivl_29123;
  tmp_ivl_29130 <= tmp_ivl_29134(1);
  tmp_ivl_29132 <= tmp_ivl_29134(0);
  tmp_ivl_29134 <= LPM_d0_ivl_29138(0 + 1 downto 0);
  tmp_ivl_29139 <= new_AGEMA_signal_2803 & n3249;
  LPM_q_ivl_29142 <= tmp_ivl_29144 & tmp_ivl_29139;
  tmp_ivl_29147 <= z2(50);
  tmp_ivl_29148 <= new_AGEMA_signal_3195 & tmp_ivl_29147;
  LPM_q_ivl_29151 <= tmp_ivl_29153 & tmp_ivl_29148;
  new_AGEMA_signal_3495 <= tmp_ivl_29155(1);
  n4126 <= tmp_ivl_29155(0);
  tmp_ivl_29155 <= LPM_d0_ivl_29159(0 + 1 downto 0);
  tmp_ivl_29161 <= z3(50);
  tmp_ivl_29162 <= new_AGEMA_signal_3564 & tmp_ivl_29161;
  LPM_q_ivl_29165 <= tmp_ivl_29167 & tmp_ivl_29162;
  tmp_ivl_29170 <= state_in_s1(202);
  tmp_ivl_29172 <= state_in_s0(202);
  tmp_ivl_29173 <= tmp_ivl_29170 & tmp_ivl_29172;
  LPM_q_ivl_29176 <= tmp_ivl_29178 & tmp_ivl_29173;
  new_AGEMA_signal_3806 <= tmp_ivl_29180(1);
  n4004 <= tmp_ivl_29180(0);
  tmp_ivl_29180 <= LPM_d0_ivl_29184(0 + 1 downto 0);
  tmp_ivl_29185 <= new_AGEMA_signal_3495 & n4126;
  LPM_q_ivl_29188 <= tmp_ivl_29190 & tmp_ivl_29185;
  tmp_ivl_29192 <= new_AGEMA_signal_3806 & n4004;
  LPM_q_ivl_29195 <= tmp_ivl_29197 & tmp_ivl_29192;
  new_AGEMA_signal_4120 <= tmp_ivl_29199(1);
  n4267 <= tmp_ivl_29199(0);
  tmp_ivl_29199 <= LPM_d0_ivl_29203(0 + 1 downto 0);
  tmp_ivl_29204 <= new_AGEMA_signal_4120 & n4267;
  LPM_q_ivl_29207 <= tmp_ivl_29209 & tmp_ivl_29204;
  tmp_ivl_29211 <= new_AGEMA_signal_4113 & n4035;
  LPM_q_ivl_29214 <= tmp_ivl_29216 & tmp_ivl_29211;
  new_AGEMA_signal_4407 <= tmp_ivl_29218(1);
  n4005 <= tmp_ivl_29218(0);
  tmp_ivl_29218 <= LPM_d0_ivl_29222(0 + 1 downto 0);
  tmp_ivl_29223 <= new_AGEMA_signal_4101 & n4006;
  LPM_q_ivl_29226 <= tmp_ivl_29228 & tmp_ivl_29223;
  tmp_ivl_29230 <= new_AGEMA_signal_4407 & n4005;
  LPM_q_ivl_29233 <= tmp_ivl_29235 & tmp_ivl_29230;
  tmp_ivl_29237 <= tmp_ivl_29241(1);
  tmp_ivl_29239 <= tmp_ivl_29241(0);
  tmp_ivl_29241 <= LPM_d0_ivl_29245(0 + 1 downto 0);
  tmp_ivl_29246 <= new_AGEMA_signal_4114 & n4046;
  LPM_q_ivl_29249 <= tmp_ivl_29251 & tmp_ivl_29246;
  tmp_ivl_29253 <= new_AGEMA_signal_4103 & n4007;
  LPM_q_ivl_29256 <= tmp_ivl_29258 & tmp_ivl_29253;
  new_AGEMA_signal_4408 <= tmp_ivl_29260(1);
  n4009 <= tmp_ivl_29260(0);
  tmp_ivl_29260 <= LPM_d0_ivl_29264(0 + 1 downto 0);
  tmp_ivl_29265 <= new_AGEMA_signal_2805 & n3248;
  LPM_q_ivl_29268 <= tmp_ivl_29270 & tmp_ivl_29265;
  tmp_ivl_29273 <= z2(51);
  tmp_ivl_29274 <= new_AGEMA_signal_3194 & tmp_ivl_29273;
  LPM_q_ivl_29277 <= tmp_ivl_29279 & tmp_ivl_29274;
  new_AGEMA_signal_3496 <= tmp_ivl_29281(1);
  n4125 <= tmp_ivl_29281(0);
  tmp_ivl_29281 <= LPM_d0_ivl_29285(0 + 1 downto 0);
  tmp_ivl_29287 <= z3(51);
  tmp_ivl_29288 <= new_AGEMA_signal_3565 & tmp_ivl_29287;
  LPM_q_ivl_29291 <= tmp_ivl_29293 & tmp_ivl_29288;
  tmp_ivl_29296 <= state_in_s1(203);
  tmp_ivl_29298 <= state_in_s0(203);
  tmp_ivl_29299 <= tmp_ivl_29296 & tmp_ivl_29298;
  LPM_q_ivl_29302 <= tmp_ivl_29304 & tmp_ivl_29299;
  new_AGEMA_signal_3807 <= tmp_ivl_29306(1);
  n4008 <= tmp_ivl_29306(0);
  tmp_ivl_29306 <= LPM_d0_ivl_29310(0 + 1 downto 0);
  tmp_ivl_29311 <= new_AGEMA_signal_3496 & n4125;
  LPM_q_ivl_29314 <= tmp_ivl_29316 & tmp_ivl_29311;
  tmp_ivl_29318 <= new_AGEMA_signal_3807 & n4008;
  LPM_q_ivl_29321 <= tmp_ivl_29323 & tmp_ivl_29318;
  new_AGEMA_signal_4121 <= tmp_ivl_29325(1);
  n4251 <= tmp_ivl_29325(0);
  tmp_ivl_29325 <= LPM_d0_ivl_29329(0 + 1 downto 0);
  tmp_ivl_29330 <= new_AGEMA_signal_4408 & n4009;
  LPM_q_ivl_29333 <= tmp_ivl_29335 & tmp_ivl_29330;
  tmp_ivl_29337 <= new_AGEMA_signal_4121 & n4251;
  LPM_q_ivl_29340 <= tmp_ivl_29342 & tmp_ivl_29337;
  tmp_ivl_29344 <= tmp_ivl_29348(1);
  tmp_ivl_29346 <= tmp_ivl_29348(0);
  tmp_ivl_29348 <= LPM_d0_ivl_29352(0 + 1 downto 0);
  tmp_ivl_29353 <= new_AGEMA_signal_4105 & n4010;
  LPM_q_ivl_29356 <= tmp_ivl_29358 & tmp_ivl_29353;
  tmp_ivl_29360 <= new_AGEMA_signal_4115 & n4050;
  LPM_q_ivl_29363 <= tmp_ivl_29365 & tmp_ivl_29360;
  new_AGEMA_signal_4409 <= tmp_ivl_29367(1);
  n4012 <= tmp_ivl_29367(0);
  tmp_ivl_29367 <= LPM_d0_ivl_29371(0 + 1 downto 0);
  tmp_ivl_29372 <= new_AGEMA_signal_2807 & n3247;
  LPM_q_ivl_29375 <= tmp_ivl_29377 & tmp_ivl_29372;
  tmp_ivl_29380 <= z2(52);
  tmp_ivl_29381 <= new_AGEMA_signal_3192 & tmp_ivl_29380;
  LPM_q_ivl_29384 <= tmp_ivl_29386 & tmp_ivl_29381;
  new_AGEMA_signal_3497 <= tmp_ivl_29388(1);
  n4123 <= tmp_ivl_29388(0);
  tmp_ivl_29388 <= LPM_d0_ivl_29392(0 + 1 downto 0);
  tmp_ivl_29394 <= z3(52);
  tmp_ivl_29395 <= new_AGEMA_signal_3566 & tmp_ivl_29394;
  LPM_q_ivl_29398 <= tmp_ivl_29400 & tmp_ivl_29395;
  tmp_ivl_29403 <= state_in_s1(204);
  tmp_ivl_29405 <= state_in_s0(204);
  tmp_ivl_29406 <= tmp_ivl_29403 & tmp_ivl_29405;
  LPM_q_ivl_29409 <= tmp_ivl_29411 & tmp_ivl_29406;
  new_AGEMA_signal_3808 <= tmp_ivl_29413(1);
  n4011 <= tmp_ivl_29413(0);
  tmp_ivl_29413 <= LPM_d0_ivl_29417(0 + 1 downto 0);
  tmp_ivl_29418 <= new_AGEMA_signal_3497 & n4123;
  LPM_q_ivl_29421 <= tmp_ivl_29423 & tmp_ivl_29418;
  tmp_ivl_29425 <= new_AGEMA_signal_3808 & n4011;
  LPM_q_ivl_29428 <= tmp_ivl_29430 & tmp_ivl_29425;
  new_AGEMA_signal_4122 <= tmp_ivl_29432(1);
  n4243 <= tmp_ivl_29432(0);
  tmp_ivl_29432 <= LPM_d0_ivl_29436(0 + 1 downto 0);
  tmp_ivl_29437 <= new_AGEMA_signal_4409 & n4012;
  LPM_q_ivl_29440 <= tmp_ivl_29442 & tmp_ivl_29437;
  tmp_ivl_29444 <= new_AGEMA_signal_4122 & n4243;
  LPM_q_ivl_29447 <= tmp_ivl_29449 & tmp_ivl_29444;
  tmp_ivl_29451 <= tmp_ivl_29455(1);
  tmp_ivl_29453 <= tmp_ivl_29455(0);
  tmp_ivl_29455 <= LPM_d0_ivl_29459(0 + 1 downto 0);
  tmp_ivl_29460 <= new_AGEMA_signal_2810 & n3246;
  LPM_q_ivl_29463 <= tmp_ivl_29465 & tmp_ivl_29460;
  tmp_ivl_29468 <= z2(53);
  tmp_ivl_29469 <= new_AGEMA_signal_3190 & tmp_ivl_29468;
  LPM_q_ivl_29472 <= tmp_ivl_29474 & tmp_ivl_29469;
  new_AGEMA_signal_3498 <= tmp_ivl_29476(1);
  n4120 <= tmp_ivl_29476(0);
  tmp_ivl_29476 <= LPM_d0_ivl_29480(0 + 1 downto 0);
  tmp_ivl_29482 <= z3(53);
  tmp_ivl_29483 <= new_AGEMA_signal_3567 & tmp_ivl_29482;
  LPM_q_ivl_29486 <= tmp_ivl_29488 & tmp_ivl_29483;
  tmp_ivl_29491 <= state_in_s1(205);
  tmp_ivl_29493 <= state_in_s0(205);
  tmp_ivl_29494 <= tmp_ivl_29491 & tmp_ivl_29493;
  LPM_q_ivl_29497 <= tmp_ivl_29499 & tmp_ivl_29494;
  new_AGEMA_signal_3809 <= tmp_ivl_29501(1);
  n4013 <= tmp_ivl_29501(0);
  tmp_ivl_29501 <= LPM_d0_ivl_29505(0 + 1 downto 0);
  tmp_ivl_29506 <= new_AGEMA_signal_3498 & n4120;
  LPM_q_ivl_29509 <= tmp_ivl_29511 & tmp_ivl_29506;
  tmp_ivl_29513 <= new_AGEMA_signal_3809 & n4013;
  LPM_q_ivl_29516 <= tmp_ivl_29518 & tmp_ivl_29513;
  new_AGEMA_signal_4123 <= tmp_ivl_29520(1);
  n4233 <= tmp_ivl_29520(0);
  tmp_ivl_29520 <= LPM_d0_ivl_29524(0 + 1 downto 0);
  tmp_ivl_29525 <= new_AGEMA_signal_4123 & n4233;
  LPM_q_ivl_29528 <= tmp_ivl_29530 & tmp_ivl_29525;
  tmp_ivl_29532 <= new_AGEMA_signal_4116 & n4055;
  LPM_q_ivl_29535 <= tmp_ivl_29537 & tmp_ivl_29532;
  new_AGEMA_signal_4410 <= tmp_ivl_29539(1);
  n4014 <= tmp_ivl_29539(0);
  tmp_ivl_29539 <= LPM_d0_ivl_29543(0 + 1 downto 0);
  tmp_ivl_29544 <= new_AGEMA_signal_4106 & n4015;
  LPM_q_ivl_29547 <= tmp_ivl_29549 & tmp_ivl_29544;
  tmp_ivl_29551 <= new_AGEMA_signal_4410 & n4014;
  LPM_q_ivl_29554 <= tmp_ivl_29556 & tmp_ivl_29551;
  tmp_ivl_29558 <= tmp_ivl_29562(1);
  tmp_ivl_29560 <= tmp_ivl_29562(0);
  tmp_ivl_29562 <= LPM_d0_ivl_29566(0 + 1 downto 0);
  tmp_ivl_29567 <= new_AGEMA_signal_2813 & n3245;
  LPM_q_ivl_29570 <= tmp_ivl_29572 & tmp_ivl_29567;
  tmp_ivl_29575 <= z2(54);
  tmp_ivl_29576 <= new_AGEMA_signal_3200 & tmp_ivl_29575;
  LPM_q_ivl_29579 <= tmp_ivl_29581 & tmp_ivl_29576;
  new_AGEMA_signal_3499 <= tmp_ivl_29583(1);
  n4118 <= tmp_ivl_29583(0);
  tmp_ivl_29583 <= LPM_d0_ivl_29587(0 + 1 downto 0);
  tmp_ivl_29589 <= z3(54);
  tmp_ivl_29590 <= new_AGEMA_signal_3568 & tmp_ivl_29589;
  LPM_q_ivl_29593 <= tmp_ivl_29595 & tmp_ivl_29590;
  tmp_ivl_29598 <= state_in_s1(206);
  tmp_ivl_29600 <= state_in_s0(206);
  tmp_ivl_29601 <= tmp_ivl_29598 & tmp_ivl_29600;
  LPM_q_ivl_29604 <= tmp_ivl_29606 & tmp_ivl_29601;
  new_AGEMA_signal_3810 <= tmp_ivl_29608(1);
  n4016 <= tmp_ivl_29608(0);
  tmp_ivl_29608 <= LPM_d0_ivl_29612(0 + 1 downto 0);
  tmp_ivl_29613 <= new_AGEMA_signal_3499 & n4118;
  LPM_q_ivl_29616 <= tmp_ivl_29618 & tmp_ivl_29613;
  tmp_ivl_29620 <= new_AGEMA_signal_3810 & n4016;
  LPM_q_ivl_29623 <= tmp_ivl_29625 & tmp_ivl_29620;
  new_AGEMA_signal_4124 <= tmp_ivl_29627(1);
  n4091 <= tmp_ivl_29627(0);
  tmp_ivl_29627 <= LPM_d0_ivl_29631(0 + 1 downto 0);
  tmp_ivl_29632 <= new_AGEMA_signal_4124 & n4091;
  LPM_q_ivl_29635 <= tmp_ivl_29637 & tmp_ivl_29632;
  tmp_ivl_29639 <= new_AGEMA_signal_4117 & n4038;
  LPM_q_ivl_29642 <= tmp_ivl_29644 & tmp_ivl_29639;
  new_AGEMA_signal_4411 <= tmp_ivl_29646(1);
  n4017 <= tmp_ivl_29646(0);
  tmp_ivl_29646 <= LPM_d0_ivl_29650(0 + 1 downto 0);
  tmp_ivl_29651 <= new_AGEMA_signal_4107 & n4018;
  LPM_q_ivl_29654 <= tmp_ivl_29656 & tmp_ivl_29651;
  tmp_ivl_29658 <= new_AGEMA_signal_4411 & n4017;
  LPM_q_ivl_29661 <= tmp_ivl_29663 & tmp_ivl_29658;
  tmp_ivl_29665 <= tmp_ivl_29669(1);
  tmp_ivl_29667 <= tmp_ivl_29669(0);
  tmp_ivl_29669 <= LPM_d0_ivl_29673(0 + 1 downto 0);
  tmp_ivl_29674 <= new_AGEMA_signal_4108 & n4019;
  LPM_q_ivl_29677 <= tmp_ivl_29679 & tmp_ivl_29674;
  tmp_ivl_29681 <= new_AGEMA_signal_4118 & n4058;
  LPM_q_ivl_29684 <= tmp_ivl_29686 & tmp_ivl_29681;
  new_AGEMA_signal_4412 <= tmp_ivl_29688(1);
  n4021 <= tmp_ivl_29688(0);
  tmp_ivl_29688 <= LPM_d0_ivl_29692(0 + 1 downto 0);
  tmp_ivl_29693 <= new_AGEMA_signal_2816 & n3244;
  LPM_q_ivl_29696 <= tmp_ivl_29698 & tmp_ivl_29693;
  tmp_ivl_29701 <= z2(55);
  tmp_ivl_29702 <= new_AGEMA_signal_3197 & tmp_ivl_29701;
  LPM_q_ivl_29705 <= tmp_ivl_29707 & tmp_ivl_29702;
  new_AGEMA_signal_3500 <= tmp_ivl_29709(1);
  n4117 <= tmp_ivl_29709(0);
  tmp_ivl_29709 <= LPM_d0_ivl_29713(0 + 1 downto 0);
  tmp_ivl_29715 <= z3(55);
  tmp_ivl_29716 <= new_AGEMA_signal_3569 & tmp_ivl_29715;
  LPM_q_ivl_29719 <= tmp_ivl_29721 & tmp_ivl_29716;
  tmp_ivl_29724 <= state_in_s1(207);
  tmp_ivl_29726 <= state_in_s0(207);
  tmp_ivl_29727 <= tmp_ivl_29724 & tmp_ivl_29726;
  LPM_q_ivl_29730 <= tmp_ivl_29732 & tmp_ivl_29727;
  new_AGEMA_signal_3811 <= tmp_ivl_29734(1);
  n4020 <= tmp_ivl_29734(0);
  tmp_ivl_29734 <= LPM_d0_ivl_29738(0 + 1 downto 0);
  tmp_ivl_29739 <= new_AGEMA_signal_3500 & n4117;
  LPM_q_ivl_29742 <= tmp_ivl_29744 & tmp_ivl_29739;
  tmp_ivl_29746 <= new_AGEMA_signal_3811 & n4020;
  LPM_q_ivl_29749 <= tmp_ivl_29751 & tmp_ivl_29746;
  new_AGEMA_signal_4125 <= tmp_ivl_29753(1);
  n4060 <= tmp_ivl_29753(0);
  tmp_ivl_29753 <= LPM_d0_ivl_29757(0 + 1 downto 0);
  tmp_ivl_29758 <= new_AGEMA_signal_4412 & n4021;
  LPM_q_ivl_29761 <= tmp_ivl_29763 & tmp_ivl_29758;
  tmp_ivl_29765 <= new_AGEMA_signal_4125 & n4060;
  LPM_q_ivl_29768 <= tmp_ivl_29770 & tmp_ivl_29765;
  tmp_ivl_29772 <= tmp_ivl_29776(1);
  tmp_ivl_29774 <= tmp_ivl_29776(0);
  tmp_ivl_29776 <= LPM_d0_ivl_29780(0 + 1 downto 0);
  tmp_ivl_29781 <= new_AGEMA_signal_2819 & n3243;
  LPM_q_ivl_29784 <= tmp_ivl_29786 & tmp_ivl_29781;
  tmp_ivl_29789 <= z2(56);
  tmp_ivl_29790 <= new_AGEMA_signal_3199 & tmp_ivl_29789;
  LPM_q_ivl_29793 <= tmp_ivl_29795 & tmp_ivl_29790;
  new_AGEMA_signal_3501 <= tmp_ivl_29797(1);
  n4114 <= tmp_ivl_29797(0);
  tmp_ivl_29797 <= LPM_d0_ivl_29801(0 + 1 downto 0);
  tmp_ivl_29803 <= z3(56);
  tmp_ivl_29804 <= new_AGEMA_signal_3570 & tmp_ivl_29803;
  LPM_q_ivl_29807 <= tmp_ivl_29809 & tmp_ivl_29804;
  tmp_ivl_29812 <= state_in_s1(192);
  tmp_ivl_29814 <= state_in_s0(192);
  tmp_ivl_29815 <= tmp_ivl_29812 & tmp_ivl_29814;
  LPM_q_ivl_29818 <= tmp_ivl_29820 & tmp_ivl_29815;
  new_AGEMA_signal_3812 <= tmp_ivl_29822(1);
  n4022 <= tmp_ivl_29822(0);
  tmp_ivl_29822 <= LPM_d0_ivl_29826(0 + 1 downto 0);
  tmp_ivl_29827 <= new_AGEMA_signal_3501 & n4114;
  LPM_q_ivl_29830 <= tmp_ivl_29832 & tmp_ivl_29827;
  tmp_ivl_29834 <= new_AGEMA_signal_3812 & n4022;
  LPM_q_ivl_29837 <= tmp_ivl_29839 & tmp_ivl_29834;
  new_AGEMA_signal_4126 <= tmp_ivl_29841(1);
  n4071 <= tmp_ivl_29841(0);
  tmp_ivl_29841 <= LPM_d0_ivl_29845(0 + 1 downto 0);
  tmp_ivl_29846 <= new_AGEMA_signal_4109 & n4023;
  LPM_q_ivl_29849 <= tmp_ivl_29851 & tmp_ivl_29846;
  tmp_ivl_29853 <= new_AGEMA_signal_4126 & n4071;
  LPM_q_ivl_29856 <= tmp_ivl_29858 & tmp_ivl_29853;
  new_AGEMA_signal_4413 <= tmp_ivl_29860(1);
  n4024 <= tmp_ivl_29860(0);
  tmp_ivl_29860 <= LPM_d0_ivl_29864(0 + 1 downto 0);
  tmp_ivl_29865 <= new_AGEMA_signal_4413 & n4024;
  LPM_q_ivl_29868 <= tmp_ivl_29870 & tmp_ivl_29865;
  tmp_ivl_29872 <= new_AGEMA_signal_4119 & n4074;
  LPM_q_ivl_29875 <= tmp_ivl_29877 & tmp_ivl_29872;
  tmp_ivl_29879 <= tmp_ivl_29883(1);
  tmp_ivl_29881 <= tmp_ivl_29883(0);
  tmp_ivl_29883 <= LPM_d0_ivl_29887(0 + 1 downto 0);
  tmp_ivl_29888 <= new_AGEMA_signal_2821 & n3242;
  LPM_q_ivl_29891 <= tmp_ivl_29893 & tmp_ivl_29888;
  tmp_ivl_29896 <= z2(57);
  tmp_ivl_29897 <= new_AGEMA_signal_3204 & tmp_ivl_29896;
  LPM_q_ivl_29900 <= tmp_ivl_29902 & tmp_ivl_29897;
  new_AGEMA_signal_3502 <= tmp_ivl_29904(1);
  n4112 <= tmp_ivl_29904(0);
  tmp_ivl_29904 <= LPM_d0_ivl_29908(0 + 1 downto 0);
  tmp_ivl_29910 <= z3(57);
  tmp_ivl_29911 <= new_AGEMA_signal_3571 & tmp_ivl_29910;
  LPM_q_ivl_29914 <= tmp_ivl_29916 & tmp_ivl_29911;
  tmp_ivl_29919 <= state_in_s1(193);
  tmp_ivl_29921 <= state_in_s0(193);
  tmp_ivl_29922 <= tmp_ivl_29919 & tmp_ivl_29921;
  LPM_q_ivl_29925 <= tmp_ivl_29927 & tmp_ivl_29922;
  new_AGEMA_signal_3813 <= tmp_ivl_29929(1);
  n4025 <= tmp_ivl_29929(0);
  tmp_ivl_29929 <= LPM_d0_ivl_29933(0 + 1 downto 0);
  tmp_ivl_29934 <= new_AGEMA_signal_3502 & n4112;
  LPM_q_ivl_29937 <= tmp_ivl_29939 & tmp_ivl_29934;
  tmp_ivl_29941 <= new_AGEMA_signal_3813 & n4025;
  LPM_q_ivl_29944 <= tmp_ivl_29946 & tmp_ivl_29941;
  new_AGEMA_signal_4127 <= tmp_ivl_29948(1);
  n4270 <= tmp_ivl_29948(0);
  tmp_ivl_29948 <= LPM_d0_ivl_29952(0 + 1 downto 0);
  tmp_ivl_29953 <= new_AGEMA_signal_4120 & n4267;
  LPM_q_ivl_29956 <= tmp_ivl_29958 & tmp_ivl_29953;
  tmp_ivl_29960 <= new_AGEMA_signal_4127 & n4270;
  LPM_q_ivl_29963 <= tmp_ivl_29965 & tmp_ivl_29960;
  new_AGEMA_signal_4414 <= tmp_ivl_29967(1);
  n4026 <= tmp_ivl_29967(0);
  tmp_ivl_29967 <= LPM_d0_ivl_29971(0 + 1 downto 0);
  tmp_ivl_29972 <= new_AGEMA_signal_4110 & n4027;
  LPM_q_ivl_29975 <= tmp_ivl_29977 & tmp_ivl_29972;
  tmp_ivl_29979 <= new_AGEMA_signal_4414 & n4026;
  LPM_q_ivl_29982 <= tmp_ivl_29984 & tmp_ivl_29979;
  tmp_ivl_29986 <= tmp_ivl_29990(1);
  tmp_ivl_29988 <= tmp_ivl_29990(0);
  tmp_ivl_29990 <= LPM_d0_ivl_29994(0 + 1 downto 0);
  tmp_ivl_29995 <= new_AGEMA_signal_2823 & n3241;
  LPM_q_ivl_29998 <= tmp_ivl_30000 & tmp_ivl_29995;
  tmp_ivl_30003 <= z2(58);
  tmp_ivl_30004 <= new_AGEMA_signal_3203 & tmp_ivl_30003;
  LPM_q_ivl_30007 <= tmp_ivl_30009 & tmp_ivl_30004;
  new_AGEMA_signal_3503 <= tmp_ivl_30011(1);
  n4226 <= tmp_ivl_30011(0);
  tmp_ivl_30011 <= LPM_d0_ivl_30015(0 + 1 downto 0);
  tmp_ivl_30017 <= z3(58);
  tmp_ivl_30018 <= new_AGEMA_signal_3572 & tmp_ivl_30017;
  LPM_q_ivl_30021 <= tmp_ivl_30023 & tmp_ivl_30018;
  tmp_ivl_30026 <= state_in_s1(194);
  tmp_ivl_30028 <= state_in_s0(194);
  tmp_ivl_30029 <= tmp_ivl_30026 & tmp_ivl_30028;
  LPM_q_ivl_30032 <= tmp_ivl_30034 & tmp_ivl_30029;
  new_AGEMA_signal_3814 <= tmp_ivl_30036(1);
  n4028 <= tmp_ivl_30036(0);
  tmp_ivl_30036 <= LPM_d0_ivl_30040(0 + 1 downto 0);
  tmp_ivl_30041 <= new_AGEMA_signal_3503 & n4226;
  LPM_q_ivl_30044 <= tmp_ivl_30046 & tmp_ivl_30041;
  tmp_ivl_30048 <= new_AGEMA_signal_3814 & n4028;
  LPM_q_ivl_30051 <= tmp_ivl_30053 & tmp_ivl_30048;
  new_AGEMA_signal_4128 <= tmp_ivl_30055(1);
  n4257 <= tmp_ivl_30055(0);
  tmp_ivl_30055 <= LPM_d0_ivl_30059(0 + 1 downto 0);
  tmp_ivl_30060 <= new_AGEMA_signal_4128 & n4257;
  LPM_q_ivl_30063 <= tmp_ivl_30065 & tmp_ivl_30060;
  tmp_ivl_30067 <= new_AGEMA_signal_4111 & n4029;
  LPM_q_ivl_30070 <= tmp_ivl_30072 & tmp_ivl_30067;
  new_AGEMA_signal_4415 <= tmp_ivl_30074(1);
  n4030 <= tmp_ivl_30074(0);
  tmp_ivl_30074 <= LPM_d0_ivl_30078(0 + 1 downto 0);
  tmp_ivl_30079 <= new_AGEMA_signal_4415 & n4030;
  LPM_q_ivl_30082 <= tmp_ivl_30084 & tmp_ivl_30079;
  tmp_ivl_30086 <= new_AGEMA_signal_4121 & n4251;
  LPM_q_ivl_30089 <= tmp_ivl_30091 & tmp_ivl_30086;
  tmp_ivl_30093 <= tmp_ivl_30097(1);
  tmp_ivl_30095 <= tmp_ivl_30097(0);
  tmp_ivl_30097 <= LPM_d0_ivl_30101(0 + 1 downto 0);
  tmp_ivl_30102 <= new_AGEMA_signal_2825 & n3240;
  LPM_q_ivl_30105 <= tmp_ivl_30107 & tmp_ivl_30102;
  tmp_ivl_30110 <= z2(59);
  tmp_ivl_30111 <= new_AGEMA_signal_3202 & tmp_ivl_30110;
  LPM_q_ivl_30114 <= tmp_ivl_30116 & tmp_ivl_30111;
  new_AGEMA_signal_3504 <= tmp_ivl_30118(1);
  n4223 <= tmp_ivl_30118(0);
  tmp_ivl_30118 <= LPM_d0_ivl_30122(0 + 1 downto 0);
  tmp_ivl_30124 <= z3(59);
  tmp_ivl_30125 <= new_AGEMA_signal_3573 & tmp_ivl_30124;
  LPM_q_ivl_30128 <= tmp_ivl_30130 & tmp_ivl_30125;
  tmp_ivl_30133 <= state_in_s1(195);
  tmp_ivl_30135 <= state_in_s0(195);
  tmp_ivl_30136 <= tmp_ivl_30133 & tmp_ivl_30135;
  LPM_q_ivl_30139 <= tmp_ivl_30141 & tmp_ivl_30136;
  new_AGEMA_signal_3815 <= tmp_ivl_30143(1);
  n4031 <= tmp_ivl_30143(0);
  tmp_ivl_30143 <= LPM_d0_ivl_30147(0 + 1 downto 0);
  tmp_ivl_30148 <= new_AGEMA_signal_3504 & n4223;
  LPM_q_ivl_30151 <= tmp_ivl_30153 & tmp_ivl_30148;
  tmp_ivl_30155 <= new_AGEMA_signal_3815 & n4031;
  LPM_q_ivl_30158 <= tmp_ivl_30160 & tmp_ivl_30155;
  new_AGEMA_signal_4129 <= tmp_ivl_30162(1);
  n4246 <= tmp_ivl_30162(0);
  tmp_ivl_30162 <= LPM_d0_ivl_30166(0 + 1 downto 0);
  tmp_ivl_30167 <= new_AGEMA_signal_4129 & n4246;
  LPM_q_ivl_30170 <= tmp_ivl_30172 & tmp_ivl_30167;
  tmp_ivl_30174 <= new_AGEMA_signal_4112 & n4032;
  LPM_q_ivl_30177 <= tmp_ivl_30179 & tmp_ivl_30174;
  new_AGEMA_signal_4416 <= tmp_ivl_30181(1);
  n4033 <= tmp_ivl_30181(0);
  tmp_ivl_30181 <= LPM_d0_ivl_30185(0 + 1 downto 0);
  tmp_ivl_30186 <= new_AGEMA_signal_4416 & n4033;
  LPM_q_ivl_30189 <= tmp_ivl_30191 & tmp_ivl_30186;
  tmp_ivl_30193 <= new_AGEMA_signal_4122 & n4243;
  LPM_q_ivl_30196 <= tmp_ivl_30198 & tmp_ivl_30193;
  tmp_ivl_30200 <= tmp_ivl_30204(1);
  tmp_ivl_30202 <= tmp_ivl_30204(0);
  tmp_ivl_30204 <= LPM_d0_ivl_30208(0 + 1 downto 0);
  tmp_ivl_30209 <= new_AGEMA_signal_2828 & n3238;
  LPM_q_ivl_30212 <= tmp_ivl_30214 & tmp_ivl_30209;
  tmp_ivl_30217 <= z2(60);
  tmp_ivl_30218 <= new_AGEMA_signal_3201 & tmp_ivl_30217;
  LPM_q_ivl_30221 <= tmp_ivl_30223 & tmp_ivl_30218;
  new_AGEMA_signal_3505 <= tmp_ivl_30225(1);
  n4220 <= tmp_ivl_30225(0);
  tmp_ivl_30225 <= LPM_d0_ivl_30229(0 + 1 downto 0);
  tmp_ivl_30231 <= z3(60);
  tmp_ivl_30232 <= new_AGEMA_signal_3575 & tmp_ivl_30231;
  LPM_q_ivl_30235 <= tmp_ivl_30237 & tmp_ivl_30232;
  tmp_ivl_30240 <= state_in_s1(196);
  tmp_ivl_30242 <= state_in_s0(196);
  tmp_ivl_30243 <= tmp_ivl_30240 & tmp_ivl_30242;
  LPM_q_ivl_30246 <= tmp_ivl_30248 & tmp_ivl_30243;
  new_AGEMA_signal_3816 <= tmp_ivl_30250(1);
  n4034 <= tmp_ivl_30250(0);
  tmp_ivl_30250 <= LPM_d0_ivl_30254(0 + 1 downto 0);
  tmp_ivl_30255 <= new_AGEMA_signal_3505 & n4220;
  LPM_q_ivl_30258 <= tmp_ivl_30260 & tmp_ivl_30255;
  tmp_ivl_30262 <= new_AGEMA_signal_3816 & n4034;
  LPM_q_ivl_30265 <= tmp_ivl_30267 & tmp_ivl_30262;
  new_AGEMA_signal_4130 <= tmp_ivl_30269(1);
  n4266 <= tmp_ivl_30269(0);
  tmp_ivl_30269 <= LPM_d0_ivl_30273(0 + 1 downto 0);
  tmp_ivl_30274 <= new_AGEMA_signal_4123 & n4233;
  LPM_q_ivl_30277 <= tmp_ivl_30279 & tmp_ivl_30274;
  tmp_ivl_30281 <= new_AGEMA_signal_4113 & n4035;
  LPM_q_ivl_30284 <= tmp_ivl_30286 & tmp_ivl_30281;
  new_AGEMA_signal_4417 <= tmp_ivl_30288(1);
  n4036 <= tmp_ivl_30288(0);
  tmp_ivl_30288 <= LPM_d0_ivl_30292(0 + 1 downto 0);
  tmp_ivl_30293 <= new_AGEMA_signal_4130 & n4266;
  LPM_q_ivl_30296 <= tmp_ivl_30298 & tmp_ivl_30293;
  tmp_ivl_30300 <= new_AGEMA_signal_4417 & n4036;
  LPM_q_ivl_30303 <= tmp_ivl_30305 & tmp_ivl_30300;
  tmp_ivl_30307 <= tmp_ivl_30311(1);
  tmp_ivl_30309 <= tmp_ivl_30311(0);
  tmp_ivl_30311 <= LPM_d0_ivl_30315(0 + 1 downto 0);
  tmp_ivl_30317 <= z2(0);
  tmp_ivl_30318 <= new_AGEMA_signal_3206 & tmp_ivl_30317;
  LPM_q_ivl_30321 <= tmp_ivl_30323 & tmp_ivl_30318;
  tmp_ivl_30325 <= new_AGEMA_signal_2831 & n4041;
  LPM_q_ivl_30328 <= tmp_ivl_30330 & tmp_ivl_30325;
  new_AGEMA_signal_3506 <= tmp_ivl_30332(1);
  n4099 <= tmp_ivl_30332(0);
  tmp_ivl_30332 <= LPM_d0_ivl_30336(0 + 1 downto 0);
  tmp_ivl_30340 <= rcon(0);
  tmp_ivl_30341 <= tmp_ivl_30337 & tmp_ivl_30340;
  LPM_q_ivl_30344 <= tmp_ivl_30346 & tmp_ivl_30341;
  tmp_ivl_30348 <= new_AGEMA_signal_3506 & n4099;
  LPM_q_ivl_30351 <= tmp_ivl_30353 & tmp_ivl_30348;
  new_AGEMA_signal_3817 <= tmp_ivl_30355(1);
  n4224 <= tmp_ivl_30355(0);
  tmp_ivl_30355 <= LPM_d0_ivl_30359(0 + 1 downto 0);
  tmp_ivl_30360 <= new_AGEMA_signal_3817 & n4224;
  LPM_q_ivl_30363 <= tmp_ivl_30365 & tmp_ivl_30360;
  tmp_ivl_30368 <= z3(0);
  tmp_ivl_30369 <= new_AGEMA_signal_3519 & tmp_ivl_30368;
  LPM_q_ivl_30372 <= tmp_ivl_30374 & tmp_ivl_30369;
  new_AGEMA_signal_4131 <= tmp_ivl_30376(1);
  n4037 <= tmp_ivl_30376(0);
  tmp_ivl_30376 <= LPM_d0_ivl_30380(0 + 1 downto 0);
  tmp_ivl_30381 <= new_AGEMA_signal_4131 & n4037;
  LPM_q_ivl_30384 <= tmp_ivl_30386 & tmp_ivl_30381;
  tmp_ivl_30389 <= state_in_s1(248);
  tmp_ivl_30391 <= state_in_s0(248);
  tmp_ivl_30392 <= tmp_ivl_30389 & tmp_ivl_30391;
  LPM_q_ivl_30395 <= tmp_ivl_30397 & tmp_ivl_30392;
  new_AGEMA_signal_4418 <= tmp_ivl_30399(1);
  n4092 <= tmp_ivl_30399(0);
  tmp_ivl_30399 <= LPM_d0_ivl_30403(0 + 1 downto 0);
  tmp_ivl_30404 <= new_AGEMA_signal_4418 & n4092;
  LPM_q_ivl_30407 <= tmp_ivl_30409 & tmp_ivl_30404;
  tmp_ivl_30411 <= new_AGEMA_signal_4127 & n4270;
  LPM_q_ivl_30414 <= tmp_ivl_30416 & tmp_ivl_30411;
  new_AGEMA_signal_4550 <= tmp_ivl_30418(1);
  n4039 <= tmp_ivl_30418(0);
  tmp_ivl_30418 <= LPM_d0_ivl_30422(0 + 1 downto 0);
  tmp_ivl_30423 <= new_AGEMA_signal_4550 & n4039;
  LPM_q_ivl_30426 <= tmp_ivl_30428 & tmp_ivl_30423;
  tmp_ivl_30430 <= new_AGEMA_signal_4117 & n4038;
  LPM_q_ivl_30433 <= tmp_ivl_30435 & tmp_ivl_30430;
  tmp_ivl_30437 <= tmp_ivl_30441(1);
  tmp_ivl_30439 <= tmp_ivl_30441(0);
  tmp_ivl_30441 <= LPM_d0_ivl_30445(0 + 1 downto 0);
  tmp_ivl_30446 <= new_AGEMA_signal_4418 & n4092;
  LPM_q_ivl_30449 <= tmp_ivl_30451 & tmp_ivl_30446;
  tmp_ivl_30453 <= new_AGEMA_signal_4102 & n4095;
  LPM_q_ivl_30456 <= tmp_ivl_30458 & tmp_ivl_30453;
  new_AGEMA_signal_4551 <= tmp_ivl_30460(1);
  n4040 <= tmp_ivl_30460(0);
  tmp_ivl_30460 <= LPM_d0_ivl_30464(0 + 1 downto 0);
  tmp_ivl_30465 <= new_AGEMA_signal_4083 & n4269;
  LPM_q_ivl_30468 <= tmp_ivl_30470 & tmp_ivl_30465;
  tmp_ivl_30472 <= new_AGEMA_signal_4551 & n4040;
  LPM_q_ivl_30475 <= tmp_ivl_30477 & tmp_ivl_30472;
  tmp_ivl_30479 <= tmp_ivl_30483(1);
  tmp_ivl_30481 <= tmp_ivl_30483(0);
  tmp_ivl_30483 <= LPM_d0_ivl_30487(0 + 1 downto 0);
  tmp_ivl_30488 <= new_AGEMA_signal_2834 & n3237;
  LPM_q_ivl_30491 <= tmp_ivl_30493 & tmp_ivl_30488;
  tmp_ivl_30496 <= z2(8);
  tmp_ivl_30497 <= new_AGEMA_signal_3294 & tmp_ivl_30496;
  LPM_q_ivl_30500 <= tmp_ivl_30502 & tmp_ivl_30497;
  new_AGEMA_signal_3507 <= tmp_ivl_30504(1);
  n4202 <= tmp_ivl_30504(0);
  tmp_ivl_30504 <= LPM_d0_ivl_30508(0 + 1 downto 0);
  tmp_ivl_30510 <= z3(8);
  tmp_ivl_30511 <= new_AGEMA_signal_3581 & tmp_ivl_30510;
  LPM_q_ivl_30514 <= tmp_ivl_30516 & tmp_ivl_30511;
  tmp_ivl_30519 <= state_in_s1(240);
  tmp_ivl_30521 <= state_in_s0(240);
  tmp_ivl_30522 <= tmp_ivl_30519 & tmp_ivl_30521;
  LPM_q_ivl_30525 <= tmp_ivl_30527 & tmp_ivl_30522;
  new_AGEMA_signal_3818 <= tmp_ivl_30529(1);
  n4042 <= tmp_ivl_30529(0);
  tmp_ivl_30529 <= LPM_d0_ivl_30533(0 + 1 downto 0);
  tmp_ivl_30534 <= new_AGEMA_signal_3507 & n4202;
  LPM_q_ivl_30537 <= tmp_ivl_30539 & tmp_ivl_30534;
  tmp_ivl_30541 <= new_AGEMA_signal_3818 & n4042;
  LPM_q_ivl_30544 <= tmp_ivl_30546 & tmp_ivl_30541;
  new_AGEMA_signal_4132 <= tmp_ivl_30548(1);
  n4061 <= tmp_ivl_30548(0);
  tmp_ivl_30548 <= LPM_d0_ivl_30552(0 + 1 downto 0);
  tmp_ivl_30553 <= new_AGEMA_signal_4104 & n4063;
  LPM_q_ivl_30556 <= tmp_ivl_30558 & tmp_ivl_30553;
  tmp_ivl_30560 <= new_AGEMA_signal_4132 & n4061;
  LPM_q_ivl_30563 <= tmp_ivl_30565 & tmp_ivl_30560;
  new_AGEMA_signal_4419 <= tmp_ivl_30567(1);
  n4043 <= tmp_ivl_30567(0);
  tmp_ivl_30567 <= LPM_d0_ivl_30571(0 + 1 downto 0);
  tmp_ivl_30572 <= new_AGEMA_signal_4098 & n4044;
  LPM_q_ivl_30575 <= tmp_ivl_30577 & tmp_ivl_30572;
  tmp_ivl_30579 <= new_AGEMA_signal_4419 & n4043;
  LPM_q_ivl_30582 <= tmp_ivl_30584 & tmp_ivl_30579;
  tmp_ivl_30586 <= tmp_ivl_30590(1);
  tmp_ivl_30588 <= tmp_ivl_30590(0);
  tmp_ivl_30590 <= LPM_d0_ivl_30594(0 + 1 downto 0);
  tmp_ivl_30595 <= new_AGEMA_signal_2837 & n3236;
  LPM_q_ivl_30598 <= tmp_ivl_30600 & tmp_ivl_30595;
  tmp_ivl_30603 <= z2(61);
  tmp_ivl_30604 <= new_AGEMA_signal_3198 & tmp_ivl_30603;
  LPM_q_ivl_30607 <= tmp_ivl_30609 & tmp_ivl_30604;
  new_AGEMA_signal_3508 <= tmp_ivl_30611(1);
  n4215 <= tmp_ivl_30611(0);
  tmp_ivl_30611 <= LPM_d0_ivl_30615(0 + 1 downto 0);
  tmp_ivl_30617 <= z3(61);
  tmp_ivl_30618 <= new_AGEMA_signal_3576 & tmp_ivl_30617;
  LPM_q_ivl_30621 <= tmp_ivl_30623 & tmp_ivl_30618;
  tmp_ivl_30626 <= state_in_s1(197);
  tmp_ivl_30628 <= state_in_s0(197);
  tmp_ivl_30629 <= tmp_ivl_30626 & tmp_ivl_30628;
  LPM_q_ivl_30632 <= tmp_ivl_30634 & tmp_ivl_30629;
  new_AGEMA_signal_3819 <= tmp_ivl_30636(1);
  n4045 <= tmp_ivl_30636(0);
  tmp_ivl_30636 <= LPM_d0_ivl_30640(0 + 1 downto 0);
  tmp_ivl_30641 <= new_AGEMA_signal_3508 & n4215;
  LPM_q_ivl_30644 <= tmp_ivl_30646 & tmp_ivl_30641;
  tmp_ivl_30648 <= new_AGEMA_signal_3819 & n4045;
  LPM_q_ivl_30651 <= tmp_ivl_30653 & tmp_ivl_30648;
  new_AGEMA_signal_4133 <= tmp_ivl_30655(1);
  n4253 <= tmp_ivl_30655(0);
  tmp_ivl_30655 <= LPM_d0_ivl_30659(0 + 1 downto 0);
  tmp_ivl_30660 <= new_AGEMA_signal_4133 & n4253;
  LPM_q_ivl_30663 <= tmp_ivl_30665 & tmp_ivl_30660;
  tmp_ivl_30667 <= new_AGEMA_signal_4124 & n4091;
  LPM_q_ivl_30670 <= tmp_ivl_30672 & tmp_ivl_30667;
  new_AGEMA_signal_4420 <= tmp_ivl_30674(1);
  n4047 <= tmp_ivl_30674(0);
  tmp_ivl_30674 <= LPM_d0_ivl_30678(0 + 1 downto 0);
  tmp_ivl_30679 <= new_AGEMA_signal_4420 & n4047;
  LPM_q_ivl_30682 <= tmp_ivl_30684 & tmp_ivl_30679;
  tmp_ivl_30686 <= new_AGEMA_signal_4114 & n4046;
  LPM_q_ivl_30689 <= tmp_ivl_30691 & tmp_ivl_30686;
  tmp_ivl_30693 <= tmp_ivl_30697(1);
  tmp_ivl_30695 <= tmp_ivl_30697(0);
  tmp_ivl_30697 <= LPM_d0_ivl_30701(0 + 1 downto 0);
  tmp_ivl_30702 <= new_AGEMA_signal_2840 & n3235;
  LPM_q_ivl_30705 <= tmp_ivl_30707 & tmp_ivl_30702;
  tmp_ivl_30710 <= z2(62);
  tmp_ivl_30711 <= new_AGEMA_signal_3209 & tmp_ivl_30710;
  LPM_q_ivl_30714 <= tmp_ivl_30716 & tmp_ivl_30711;
  new_AGEMA_signal_3509 <= tmp_ivl_30718(1);
  n4107 <= tmp_ivl_30718(0);
  tmp_ivl_30718 <= LPM_d0_ivl_30722(0 + 1 downto 0);
  tmp_ivl_30723 <= new_AGEMA_signal_3509 & n4107;
  LPM_q_ivl_30726 <= tmp_ivl_30728 & tmp_ivl_30723;
  tmp_ivl_30731 <= z3(62);
  tmp_ivl_30732 <= new_AGEMA_signal_3577 & tmp_ivl_30731;
  LPM_q_ivl_30735 <= tmp_ivl_30737 & tmp_ivl_30732;
  new_AGEMA_signal_3820 <= tmp_ivl_30739(1);
  n4048 <= tmp_ivl_30739(0);
  tmp_ivl_30739 <= LPM_d0_ivl_30743(0 + 1 downto 0);
  tmp_ivl_30744 <= new_AGEMA_signal_3820 & n4048;
  LPM_q_ivl_30747 <= tmp_ivl_30749 & tmp_ivl_30744;
  tmp_ivl_30752 <= state_in_s1(198);
  tmp_ivl_30754 <= state_in_s0(198);
  tmp_ivl_30755 <= tmp_ivl_30752 & tmp_ivl_30754;
  LPM_q_ivl_30758 <= tmp_ivl_30760 & tmp_ivl_30755;
  new_AGEMA_signal_4134 <= tmp_ivl_30762(1);
  n4242 <= tmp_ivl_30762(0);
  tmp_ivl_30762 <= LPM_d0_ivl_30766(0 + 1 downto 0);
  tmp_ivl_30767 <= new_AGEMA_signal_4132 & n4061;
  LPM_q_ivl_30770 <= tmp_ivl_30772 & tmp_ivl_30767;
  tmp_ivl_30774 <= new_AGEMA_signal_4134 & n4242;
  LPM_q_ivl_30777 <= tmp_ivl_30779 & tmp_ivl_30774;
  new_AGEMA_signal_4421 <= tmp_ivl_30781(1);
  n4049 <= tmp_ivl_30781(0);
  tmp_ivl_30781 <= LPM_d0_ivl_30785(0 + 1 downto 0);
  tmp_ivl_30786 <= new_AGEMA_signal_4097 & n4239;
  LPM_q_ivl_30789 <= tmp_ivl_30791 & tmp_ivl_30786;
  tmp_ivl_30793 <= new_AGEMA_signal_4421 & n4049;
  LPM_q_ivl_30796 <= tmp_ivl_30798 & tmp_ivl_30793;
  tmp_ivl_30800 <= tmp_ivl_30804(1);
  tmp_ivl_30802 <= tmp_ivl_30804(0);
  tmp_ivl_30804 <= LPM_d0_ivl_30808(0 + 1 downto 0);
  tmp_ivl_30809 <= new_AGEMA_signal_4115 & n4050;
  LPM_q_ivl_30812 <= tmp_ivl_30814 & tmp_ivl_30809;
  tmp_ivl_30816 <= new_AGEMA_signal_4134 & n4242;
  LPM_q_ivl_30819 <= tmp_ivl_30821 & tmp_ivl_30816;
  new_AGEMA_signal_4422 <= tmp_ivl_30823(1);
  n4051 <= tmp_ivl_30823(0);
  tmp_ivl_30823 <= LPM_d0_ivl_30827(0 + 1 downto 0);
  tmp_ivl_30828 <= new_AGEMA_signal_4125 & n4060;
  LPM_q_ivl_30831 <= tmp_ivl_30833 & tmp_ivl_30828;
  tmp_ivl_30835 <= new_AGEMA_signal_4422 & n4051;
  LPM_q_ivl_30838 <= tmp_ivl_30840 & tmp_ivl_30835;
  tmp_ivl_30842 <= tmp_ivl_30846(1);
  tmp_ivl_30844 <= tmp_ivl_30846(0);
  tmp_ivl_30846 <= LPM_d0_ivl_30850(0 + 1 downto 0);
  tmp_ivl_30852 <= z2(4);
  tmp_ivl_30853 <= new_AGEMA_signal_3208 & tmp_ivl_30852;
  LPM_q_ivl_30856 <= tmp_ivl_30858 & tmp_ivl_30853;
  tmp_ivl_30860 <= new_AGEMA_signal_2990 & n3232;
  LPM_q_ivl_30863 <= tmp_ivl_30865 & tmp_ivl_30860;
  new_AGEMA_signal_3510 <= tmp_ivl_30867(1);
  n4250 <= tmp_ivl_30867(0);
  tmp_ivl_30867 <= LPM_d0_ivl_30871(0 + 1 downto 0);
  tmp_ivl_30872 <= new_AGEMA_signal_2846 & n3234;
  LPM_q_ivl_30875 <= tmp_ivl_30877 & tmp_ivl_30872;
  tmp_ivl_30880 <= z2(63);
  tmp_ivl_30881 <= new_AGEMA_signal_3205 & tmp_ivl_30880;
  LPM_q_ivl_30884 <= tmp_ivl_30886 & tmp_ivl_30881;
  new_AGEMA_signal_3511 <= tmp_ivl_30888(1);
  n4104 <= tmp_ivl_30888(0);
  tmp_ivl_30888 <= LPM_d0_ivl_30892(0 + 1 downto 0);
  tmp_ivl_30893 <= new_AGEMA_signal_3511 & n4104;
  LPM_q_ivl_30896 <= tmp_ivl_30898 & tmp_ivl_30893;
  tmp_ivl_30900 <= new_AGEMA_signal_3509 & n4107;
  LPM_q_ivl_30903 <= tmp_ivl_30905 & tmp_ivl_30900;
  new_AGEMA_signal_3821 <= tmp_ivl_30907(1);
  n4052 <= tmp_ivl_30907(0);
  tmp_ivl_30907 <= LPM_d0_ivl_30911(0 + 1 downto 0);
  tmp_ivl_30912 <= new_AGEMA_signal_3510 & n4250;
  LPM_q_ivl_30915 <= tmp_ivl_30917 & tmp_ivl_30912;
  tmp_ivl_30919 <= new_AGEMA_signal_3821 & n4052;
  LPM_q_ivl_30922 <= tmp_ivl_30924 & tmp_ivl_30919;
  tmp_ivl_30926 <= tmp_ivl_30930(1);
  tmp_ivl_30928 <= tmp_ivl_30930(0);
  tmp_ivl_30930 <= LPM_d0_ivl_30934(0 + 1 downto 0);
  tmp_ivl_30935 <= new_AGEMA_signal_4079 & n4072;
  LPM_q_ivl_30938 <= tmp_ivl_30940 & tmp_ivl_30935;
  tmp_ivl_30942 <= new_AGEMA_signal_4100 & n4229;
  LPM_q_ivl_30945 <= tmp_ivl_30947 & tmp_ivl_30942;
  new_AGEMA_signal_4423 <= tmp_ivl_30949(1);
  n4054 <= tmp_ivl_30949(0);
  tmp_ivl_30949 <= LPM_d0_ivl_30953(0 + 1 downto 0);
  tmp_ivl_30955 <= z3(63);
  tmp_ivl_30956 <= new_AGEMA_signal_3578 & tmp_ivl_30955;
  LPM_q_ivl_30959 <= tmp_ivl_30961 & tmp_ivl_30956;
  tmp_ivl_30964 <= state_in_s1(199);
  tmp_ivl_30966 <= state_in_s0(199);
  tmp_ivl_30967 <= tmp_ivl_30964 & tmp_ivl_30966;
  LPM_q_ivl_30970 <= tmp_ivl_30972 & tmp_ivl_30967;
  new_AGEMA_signal_3822 <= tmp_ivl_30974(1);
  n4053 <= tmp_ivl_30974(0);
  tmp_ivl_30974 <= LPM_d0_ivl_30978(0 + 1 downto 0);
  tmp_ivl_30979 <= new_AGEMA_signal_3511 & n4104;
  LPM_q_ivl_30982 <= tmp_ivl_30984 & tmp_ivl_30979;
  tmp_ivl_30986 <= new_AGEMA_signal_3822 & n4053;
  LPM_q_ivl_30989 <= tmp_ivl_30991 & tmp_ivl_30986;
  new_AGEMA_signal_4136 <= tmp_ivl_30993(1);
  n4232 <= tmp_ivl_30993(0);
  tmp_ivl_30993 <= LPM_d0_ivl_30997(0 + 1 downto 0);
  tmp_ivl_30998 <= new_AGEMA_signal_4423 & n4054;
  LPM_q_ivl_31001 <= tmp_ivl_31003 & tmp_ivl_30998;
  tmp_ivl_31005 <= new_AGEMA_signal_4136 & n4232;
  LPM_q_ivl_31008 <= tmp_ivl_31010 & tmp_ivl_31005;
  tmp_ivl_31012 <= tmp_ivl_31016(1);
  tmp_ivl_31014 <= tmp_ivl_31016(0);
  tmp_ivl_31016 <= LPM_d0_ivl_31020(0 + 1 downto 0);
  tmp_ivl_31021 <= new_AGEMA_signal_4136 & n4232;
  LPM_q_ivl_31024 <= tmp_ivl_31026 & tmp_ivl_31021;
  tmp_ivl_31028 <= new_AGEMA_signal_4116 & n4055;
  LPM_q_ivl_31031 <= tmp_ivl_31033 & tmp_ivl_31028;
  new_AGEMA_signal_4424 <= tmp_ivl_31035(1);
  n4056 <= tmp_ivl_31035(0);
  tmp_ivl_31035 <= LPM_d0_ivl_31039(0 + 1 downto 0);
  tmp_ivl_31040 <= new_AGEMA_signal_4126 & n4071;
  LPM_q_ivl_31043 <= tmp_ivl_31045 & tmp_ivl_31040;
  tmp_ivl_31047 <= new_AGEMA_signal_4424 & n4056;
  LPM_q_ivl_31050 <= tmp_ivl_31052 & tmp_ivl_31047;
  tmp_ivl_31054 <= tmp_ivl_31058(1);
  tmp_ivl_31056 <= tmp_ivl_31058(0);
  tmp_ivl_31058 <= LPM_d0_ivl_31062(0 + 1 downto 0);
  tmp_ivl_31064 <= z2(1);
  tmp_ivl_31065 <= new_AGEMA_signal_3212 & tmp_ivl_31064;
  LPM_q_ivl_31068 <= tmp_ivl_31070 & tmp_ivl_31065;
  tmp_ivl_31072 <= new_AGEMA_signal_2849 & n4066;
  LPM_q_ivl_31075 <= tmp_ivl_31077 & tmp_ivl_31072;
  new_AGEMA_signal_3512 <= tmp_ivl_31079(1);
  n4101 <= tmp_ivl_31079(0);
  tmp_ivl_31079 <= LPM_d0_ivl_31083(0 + 1 downto 0);
  tmp_ivl_31086 <= tmp_ivl_31084 & n4206;
  LPM_q_ivl_31089 <= tmp_ivl_31091 & tmp_ivl_31086;
  tmp_ivl_31093 <= new_AGEMA_signal_3512 & n4101;
  LPM_q_ivl_31096 <= tmp_ivl_31098 & tmp_ivl_31093;
  new_AGEMA_signal_3823 <= tmp_ivl_31100(1);
  n4222 <= tmp_ivl_31100(0);
  tmp_ivl_31100 <= LPM_d0_ivl_31104(0 + 1 downto 0);
  tmp_ivl_31105 <= new_AGEMA_signal_3823 & n4222;
  LPM_q_ivl_31108 <= tmp_ivl_31110 & tmp_ivl_31105;
  tmp_ivl_31113 <= z3(1);
  tmp_ivl_31114 <= new_AGEMA_signal_3530 & tmp_ivl_31113;
  LPM_q_ivl_31117 <= tmp_ivl_31119 & tmp_ivl_31114;
  new_AGEMA_signal_4137 <= tmp_ivl_31121(1);
  n4057 <= tmp_ivl_31121(0);
  tmp_ivl_31121 <= LPM_d0_ivl_31125(0 + 1 downto 0);
  tmp_ivl_31127 <= state_in_s1(249);
  tmp_ivl_31129 <= state_in_s0(249);
  tmp_ivl_31130 <= tmp_ivl_31127 & tmp_ivl_31129;
  LPM_q_ivl_31133 <= tmp_ivl_31135 & tmp_ivl_31130;
  tmp_ivl_31137 <= new_AGEMA_signal_4137 & n4057;
  LPM_q_ivl_31140 <= tmp_ivl_31142 & tmp_ivl_31137;
  new_AGEMA_signal_4425 <= tmp_ivl_31144(1);
  n4065 <= tmp_ivl_31144(0);
  tmp_ivl_31144 <= LPM_d0_ivl_31148(0 + 1 downto 0);
  tmp_ivl_31149 <= new_AGEMA_signal_4128 & n4257;
  LPM_q_ivl_31152 <= tmp_ivl_31154 & tmp_ivl_31149;
  tmp_ivl_31156 <= new_AGEMA_signal_4425 & n4065;
  LPM_q_ivl_31159 <= tmp_ivl_31161 & tmp_ivl_31156;
  new_AGEMA_signal_4558 <= tmp_ivl_31163(1);
  n4059 <= tmp_ivl_31163(0);
  tmp_ivl_31163 <= LPM_d0_ivl_31167(0 + 1 downto 0);
  tmp_ivl_31168 <= new_AGEMA_signal_4558 & n4059;
  LPM_q_ivl_31171 <= tmp_ivl_31173 & tmp_ivl_31168;
  tmp_ivl_31175 <= new_AGEMA_signal_4118 & n4058;
  LPM_q_ivl_31178 <= tmp_ivl_31180 & tmp_ivl_31175;
  tmp_ivl_31182 <= tmp_ivl_31186(1);
  tmp_ivl_31184 <= tmp_ivl_31186(0);
  tmp_ivl_31186 <= LPM_d0_ivl_31190(0 + 1 downto 0);
  tmp_ivl_31191 <= new_AGEMA_signal_4132 & n4061;
  LPM_q_ivl_31194 <= tmp_ivl_31196 & tmp_ivl_31191;
  tmp_ivl_31198 <= new_AGEMA_signal_4125 & n4060;
  LPM_q_ivl_31201 <= tmp_ivl_31203 & tmp_ivl_31198;
  new_AGEMA_signal_4426 <= tmp_ivl_31205(1);
  n4062 <= tmp_ivl_31205(0);
  tmp_ivl_31205 <= LPM_d0_ivl_31209(0 + 1 downto 0);
  tmp_ivl_31210 <= new_AGEMA_signal_4426 & n4062;
  LPM_q_ivl_31213 <= tmp_ivl_31215 & tmp_ivl_31210;
  tmp_ivl_31217 <= new_AGEMA_signal_4425 & n4065;
  LPM_q_ivl_31220 <= tmp_ivl_31222 & tmp_ivl_31217;
  tmp_ivl_31224 <= tmp_ivl_31228(1);
  tmp_ivl_31226 <= tmp_ivl_31228(0);
  tmp_ivl_31228 <= LPM_d0_ivl_31232(0 + 1 downto 0);
  tmp_ivl_31233 <= new_AGEMA_signal_4085 & n4258;
  LPM_q_ivl_31236 <= tmp_ivl_31238 & tmp_ivl_31233;
  tmp_ivl_31240 <= new_AGEMA_signal_4104 & n4063;
  LPM_q_ivl_31243 <= tmp_ivl_31245 & tmp_ivl_31240;
  new_AGEMA_signal_4427 <= tmp_ivl_31247(1);
  n4064 <= tmp_ivl_31247(0);
  tmp_ivl_31247 <= LPM_d0_ivl_31251(0 + 1 downto 0);
  tmp_ivl_31252 <= new_AGEMA_signal_4425 & n4065;
  LPM_q_ivl_31255 <= tmp_ivl_31257 & tmp_ivl_31252;
  tmp_ivl_31259 <= new_AGEMA_signal_4427 & n4064;
  LPM_q_ivl_31262 <= tmp_ivl_31264 & tmp_ivl_31259;
  tmp_ivl_31266 <= tmp_ivl_31270(1);
  tmp_ivl_31268 <= tmp_ivl_31270(0);
  tmp_ivl_31270 <= LPM_d0_ivl_31274(0 + 1 downto 0);
  tmp_ivl_31276 <= z2(2);
  tmp_ivl_31277 <= new_AGEMA_signal_3211 & tmp_ivl_31276;
  LPM_q_ivl_31280 <= tmp_ivl_31282 & tmp_ivl_31277;
  tmp_ivl_31284 <= new_AGEMA_signal_3824 & n3287;
  LPM_q_ivl_31287 <= tmp_ivl_31289 & tmp_ivl_31284;
  new_AGEMA_signal_4138 <= tmp_ivl_31291(1);
  n4217 <= tmp_ivl_31291(0);
  tmp_ivl_31291 <= LPM_d0_ivl_31295(0 + 1 downto 0);
  tmp_ivl_31297 <= z3(2);
  tmp_ivl_31298 <= new_AGEMA_signal_3541 & tmp_ivl_31297;
  LPM_q_ivl_31301 <= tmp_ivl_31303 & tmp_ivl_31298;
  tmp_ivl_31306 <= state_in_s1(250);
  tmp_ivl_31308 <= state_in_s0(250);
  tmp_ivl_31309 <= tmp_ivl_31306 & tmp_ivl_31308;
  LPM_q_ivl_31312 <= tmp_ivl_31314 & tmp_ivl_31309;
  new_AGEMA_signal_3825 <= tmp_ivl_31316(1);
  n4070 <= tmp_ivl_31316(0);
  tmp_ivl_31316 <= LPM_d0_ivl_31320(0 + 1 downto 0);
  tmp_ivl_31321 <= new_AGEMA_signal_4138 & n4217;
  LPM_q_ivl_31324 <= tmp_ivl_31326 & tmp_ivl_31321;
  tmp_ivl_31328 <= new_AGEMA_signal_3825 & n4070;
  LPM_q_ivl_31331 <= tmp_ivl_31333 & tmp_ivl_31328;
  new_AGEMA_signal_4428 <= tmp_ivl_31335(1);
  n4078 <= tmp_ivl_31335(0);
  tmp_ivl_31335 <= LPM_d0_ivl_31339(0 + 1 downto 0);
  tmp_ivl_31340 <= new_AGEMA_signal_4079 & n4072;
  LPM_q_ivl_31343 <= tmp_ivl_31345 & tmp_ivl_31340;
  tmp_ivl_31347 <= new_AGEMA_signal_4126 & n4071;
  LPM_q_ivl_31350 <= tmp_ivl_31352 & tmp_ivl_31347;
  new_AGEMA_signal_4429 <= tmp_ivl_31354(1);
  n4073 <= tmp_ivl_31354(0);
  tmp_ivl_31354 <= LPM_d0_ivl_31358(0 + 1 downto 0);
  tmp_ivl_31359 <= new_AGEMA_signal_4428 & n4078;
  LPM_q_ivl_31362 <= tmp_ivl_31364 & tmp_ivl_31359;
  tmp_ivl_31366 <= new_AGEMA_signal_4429 & n4073;
  LPM_q_ivl_31369 <= tmp_ivl_31371 & tmp_ivl_31366;
  tmp_ivl_31373 <= tmp_ivl_31377(1);
  tmp_ivl_31375 <= tmp_ivl_31377(0);
  tmp_ivl_31377 <= LPM_d0_ivl_31381(0 + 1 downto 0);
  tmp_ivl_31382 <= new_AGEMA_signal_4129 & n4246;
  LPM_q_ivl_31385 <= tmp_ivl_31387 & tmp_ivl_31382;
  tmp_ivl_31389 <= new_AGEMA_signal_4119 & n4074;
  LPM_q_ivl_31392 <= tmp_ivl_31394 & tmp_ivl_31389;
  new_AGEMA_signal_4430 <= tmp_ivl_31396(1);
  n4075 <= tmp_ivl_31396(0);
  tmp_ivl_31396 <= LPM_d0_ivl_31400(0 + 1 downto 0);
  tmp_ivl_31401 <= new_AGEMA_signal_4428 & n4078;
  LPM_q_ivl_31404 <= tmp_ivl_31406 & tmp_ivl_31401;
  tmp_ivl_31408 <= new_AGEMA_signal_4430 & n4075;
  LPM_q_ivl_31411 <= tmp_ivl_31413 & tmp_ivl_31408;
  tmp_ivl_31415 <= tmp_ivl_31419(1);
  tmp_ivl_31417 <= tmp_ivl_31419(0);
  tmp_ivl_31419 <= LPM_d0_ivl_31423(0 + 1 downto 0);
  tmp_ivl_31424 <= new_AGEMA_signal_4088 & n4245;
  LPM_q_ivl_31427 <= tmp_ivl_31429 & tmp_ivl_31424;
  tmp_ivl_31431 <= new_AGEMA_signal_4080 & n4076;
  LPM_q_ivl_31434 <= tmp_ivl_31436 & tmp_ivl_31431;
  new_AGEMA_signal_4431 <= tmp_ivl_31438(1);
  n4077 <= tmp_ivl_31438(0);
  tmp_ivl_31438 <= LPM_d0_ivl_31442(0 + 1 downto 0);
  tmp_ivl_31443 <= new_AGEMA_signal_4428 & n4078;
  LPM_q_ivl_31446 <= tmp_ivl_31448 & tmp_ivl_31443;
  tmp_ivl_31450 <= new_AGEMA_signal_4431 & n4077;
  LPM_q_ivl_31453 <= tmp_ivl_31455 & tmp_ivl_31450;
  tmp_ivl_31457 <= tmp_ivl_31461(1);
  tmp_ivl_31459 <= tmp_ivl_31461(0);
  tmp_ivl_31461 <= LPM_d0_ivl_31465(0 + 1 downto 0);
  tmp_ivl_31467 <= z2(3);
  tmp_ivl_31468 <= new_AGEMA_signal_3210 & tmp_ivl_31467;
  LPM_q_ivl_31471 <= tmp_ivl_31473 & tmp_ivl_31468;
  tmp_ivl_31475 <= new_AGEMA_signal_4432 & n3233;
  LPM_q_ivl_31478 <= tmp_ivl_31480 & tmp_ivl_31475;
  new_AGEMA_signal_4564 <= tmp_ivl_31482(1);
  n4262 <= tmp_ivl_31482(0);
  tmp_ivl_31482 <= LPM_d0_ivl_31486(0 + 1 downto 0);
  tmp_ivl_31487 <= new_AGEMA_signal_3508 & n4215;
  LPM_q_ivl_31490 <= tmp_ivl_31492 & tmp_ivl_31487;
  tmp_ivl_31494 <= new_AGEMA_signal_4564 & n4262;
  LPM_q_ivl_31497 <= tmp_ivl_31499 & tmp_ivl_31494;
  new_AGEMA_signal_4602 <= tmp_ivl_31501(1);
  n4082 <= tmp_ivl_31501(0);
  tmp_ivl_31501 <= LPM_d0_ivl_31505(0 + 1 downto 0);
  tmp_ivl_31506 <= new_AGEMA_signal_4602 & n4082;
  LPM_q_ivl_31509 <= tmp_ivl_31511 & tmp_ivl_31506;
  tmp_ivl_31513 <= new_AGEMA_signal_3509 & n4107;
  LPM_q_ivl_31516 <= tmp_ivl_31518 & tmp_ivl_31513;
  tmp_ivl_31520 <= tmp_ivl_31524(1);
  tmp_ivl_31522 <= tmp_ivl_31524(0);
  tmp_ivl_31524 <= LPM_d0_ivl_31528(0 + 1 downto 0);
  tmp_ivl_31529 <= new_AGEMA_signal_4564 & n4262;
  LPM_q_ivl_31532 <= tmp_ivl_31534 & tmp_ivl_31529;
  tmp_ivl_31536 <= new_AGEMA_signal_4138 & n4217;
  LPM_q_ivl_31539 <= tmp_ivl_31541 & tmp_ivl_31536;
  new_AGEMA_signal_4603 <= tmp_ivl_31543(1);
  n4083 <= tmp_ivl_31543(0);
  tmp_ivl_31543 <= LPM_d0_ivl_31547(0 + 1 downto 0);
  tmp_ivl_31548 <= new_AGEMA_signal_4603 & n4083;
  LPM_q_ivl_31551 <= tmp_ivl_31553 & tmp_ivl_31548;
  tmp_ivl_31555 <= new_AGEMA_signal_3507 & n4202;
  LPM_q_ivl_31558 <= tmp_ivl_31560 & tmp_ivl_31555;
  tmp_ivl_31562 <= tmp_ivl_31566(1);
  tmp_ivl_31564 <= tmp_ivl_31566(0);
  tmp_ivl_31566 <= LPM_d0_ivl_31570(0 + 1 downto 0);
  tmp_ivl_31571 <= new_AGEMA_signal_4433 & n3239;
  LPM_q_ivl_31574 <= tmp_ivl_31576 & tmp_ivl_31571;
  tmp_ivl_31579 <= z2(7);
  tmp_ivl_31580 <= new_AGEMA_signal_3269 & tmp_ivl_31579;
  LPM_q_ivl_31583 <= tmp_ivl_31585 & tmp_ivl_31580;
  new_AGEMA_signal_4565 <= tmp_ivl_31587(1);
  n4219 <= tmp_ivl_31587(0);
  tmp_ivl_31587 <= LPM_d0_ivl_31591(0 + 1 downto 0);
  tmp_ivl_31592 <= new_AGEMA_signal_4565 & n4219;
  LPM_q_ivl_31595 <= tmp_ivl_31597 & tmp_ivl_31592;
  tmp_ivl_31599 <= new_AGEMA_signal_3463 & n4192;
  LPM_q_ivl_31602 <= tmp_ivl_31604 & tmp_ivl_31599;
  new_AGEMA_signal_4604 <= tmp_ivl_31606(1);
  n4088 <= tmp_ivl_31606(0);
  tmp_ivl_31606 <= LPM_d0_ivl_31610(0 + 1 downto 0);
  tmp_ivl_31611 <= new_AGEMA_signal_3826 & n3230;
  LPM_q_ivl_31614 <= tmp_ivl_31616 & tmp_ivl_31611;
  tmp_ivl_31619 <= z2(6);
  tmp_ivl_31620 <= new_AGEMA_signal_3272 & tmp_ivl_31619;
  LPM_q_ivl_31623 <= tmp_ivl_31625 & tmp_ivl_31620;
  new_AGEMA_signal_4143 <= tmp_ivl_31627(1);
  n4228 <= tmp_ivl_31627(0);
  tmp_ivl_31627 <= LPM_d0_ivl_31631(0 + 1 downto 0);
  tmp_ivl_31632 <= new_AGEMA_signal_4604 & n4088;
  LPM_q_ivl_31635 <= tmp_ivl_31637 & tmp_ivl_31632;
  tmp_ivl_31639 <= new_AGEMA_signal_4143 & n4228;
  LPM_q_ivl_31642 <= tmp_ivl_31644 & tmp_ivl_31639;
  tmp_ivl_31646 <= tmp_ivl_31650(1);
  tmp_ivl_31648 <= tmp_ivl_31650(0);
  tmp_ivl_31650 <= LPM_d0_ivl_31654(0 + 1 downto 0);
  tmp_ivl_31656 <= z3(7);
  tmp_ivl_31657 <= new_AGEMA_signal_3580 & tmp_ivl_31656;
  LPM_q_ivl_31660 <= tmp_ivl_31662 & tmp_ivl_31657;
  tmp_ivl_31665 <= state_in_s1(255);
  tmp_ivl_31667 <= state_in_s0(255);
  tmp_ivl_31668 <= tmp_ivl_31665 & tmp_ivl_31667;
  LPM_q_ivl_31671 <= tmp_ivl_31673 & tmp_ivl_31668;
  new_AGEMA_signal_3827 <= tmp_ivl_31675(1);
  n4089 <= tmp_ivl_31675(0);
  tmp_ivl_31675 <= LPM_d0_ivl_31679(0 + 1 downto 0);
  tmp_ivl_31680 <= new_AGEMA_signal_4565 & n4219;
  LPM_q_ivl_31683 <= tmp_ivl_31685 & tmp_ivl_31680;
  tmp_ivl_31687 <= new_AGEMA_signal_3827 & n4089;
  LPM_q_ivl_31690 <= tmp_ivl_31692 & tmp_ivl_31687;
  new_AGEMA_signal_4605 <= tmp_ivl_31694(1);
  n4097 <= tmp_ivl_31694(0);
  tmp_ivl_31694 <= LPM_d0_ivl_31698(0 + 1 downto 0);
  tmp_ivl_31699 <= new_AGEMA_signal_4133 & n4253;
  LPM_q_ivl_31702 <= tmp_ivl_31704 & tmp_ivl_31699;
  tmp_ivl_31706 <= new_AGEMA_signal_4605 & n4097;
  LPM_q_ivl_31709 <= tmp_ivl_31711 & tmp_ivl_31706;
  new_AGEMA_signal_4627 <= tmp_ivl_31713(1);
  n4090 <= tmp_ivl_31713(0);
  tmp_ivl_31713 <= LPM_d0_ivl_31717(0 + 1 downto 0);
  tmp_ivl_31718 <= new_AGEMA_signal_4094 & n4255;
  LPM_q_ivl_31721 <= tmp_ivl_31723 & tmp_ivl_31718;
  tmp_ivl_31725 <= new_AGEMA_signal_4627 & n4090;
  LPM_q_ivl_31728 <= tmp_ivl_31730 & tmp_ivl_31725;
  tmp_ivl_31732 <= tmp_ivl_31736(1);
  tmp_ivl_31734 <= tmp_ivl_31736(0);
  tmp_ivl_31736 <= LPM_d0_ivl_31740(0 + 1 downto 0);
  tmp_ivl_31741 <= new_AGEMA_signal_4605 & n4097;
  LPM_q_ivl_31744 <= tmp_ivl_31746 & tmp_ivl_31741;
  tmp_ivl_31748 <= new_AGEMA_signal_4124 & n4091;
  LPM_q_ivl_31751 <= tmp_ivl_31753 & tmp_ivl_31748;
  new_AGEMA_signal_4628 <= tmp_ivl_31755(1);
  n4093 <= tmp_ivl_31755(0);
  tmp_ivl_31755 <= LPM_d0_ivl_31759(0 + 1 downto 0);
  tmp_ivl_31760 <= new_AGEMA_signal_4628 & n4093;
  LPM_q_ivl_31763 <= tmp_ivl_31765 & tmp_ivl_31760;
  tmp_ivl_31767 <= new_AGEMA_signal_4418 & n4092;
  LPM_q_ivl_31770 <= tmp_ivl_31772 & tmp_ivl_31767;
  tmp_ivl_31774 <= tmp_ivl_31778(1);
  tmp_ivl_31776 <= tmp_ivl_31778(0);
  tmp_ivl_31778 <= LPM_d0_ivl_31782(0 + 1 downto 0);
  tmp_ivl_31783 <= new_AGEMA_signal_4102 & n4095;
  LPM_q_ivl_31786 <= tmp_ivl_31788 & tmp_ivl_31783;
  tmp_ivl_31790 <= new_AGEMA_signal_4095 & n4094;
  LPM_q_ivl_31793 <= tmp_ivl_31795 & tmp_ivl_31790;
  new_AGEMA_signal_4434 <= tmp_ivl_31797(1);
  n4096 <= tmp_ivl_31797(0);
  tmp_ivl_31797 <= LPM_d0_ivl_31801(0 + 1 downto 0);
  tmp_ivl_31802 <= new_AGEMA_signal_4605 & n4097;
  LPM_q_ivl_31805 <= tmp_ivl_31807 & tmp_ivl_31802;
  tmp_ivl_31809 <= new_AGEMA_signal_4434 & n4096;
  LPM_q_ivl_31812 <= tmp_ivl_31814 & tmp_ivl_31809;
  tmp_ivl_31816 <= tmp_ivl_31820(1);
  tmp_ivl_31818 <= tmp_ivl_31820(0);
  tmp_ivl_31820 <= LPM_d0_ivl_31824(0 + 1 downto 0);
  tmp_ivl_31825 <= new_AGEMA_signal_3511 & n4104;
  LPM_q_ivl_31828 <= tmp_ivl_31830 & tmp_ivl_31825;
  tmp_ivl_31832 <= new_AGEMA_signal_3506 & n4099;
  LPM_q_ivl_31835 <= tmp_ivl_31837 & tmp_ivl_31832;
  new_AGEMA_signal_3828 <= tmp_ivl_31839(1);
  n4098 <= tmp_ivl_31839(0);
  tmp_ivl_31839 <= LPM_d0_ivl_31843(0 + 1 downto 0);
  tmp_ivl_31845 <= z2(5);
  tmp_ivl_31846 <= new_AGEMA_signal_3207 & tmp_ivl_31845;
  LPM_q_ivl_31849 <= tmp_ivl_31851 & tmp_ivl_31846;
  tmp_ivl_31853 <= new_AGEMA_signal_2858 & n4103;
  LPM_q_ivl_31856 <= tmp_ivl_31858 & tmp_ivl_31853;
  new_AGEMA_signal_3514 <= tmp_ivl_31860(1);
  n4205 <= tmp_ivl_31860(0);
  tmp_ivl_31860 <= LPM_d0_ivl_31864(0 + 1 downto 0);
  tmp_ivl_31868 <= rcon(1);
  tmp_ivl_31869 <= tmp_ivl_31865 & tmp_ivl_31868;
  LPM_q_ivl_31872 <= tmp_ivl_31874 & tmp_ivl_31869;
  tmp_ivl_31876 <= new_AGEMA_signal_3514 & n4205;
  LPM_q_ivl_31879 <= tmp_ivl_31881 & tmp_ivl_31876;
  new_AGEMA_signal_3829 <= tmp_ivl_31883(1);
  n4210 <= tmp_ivl_31883(0);
  tmp_ivl_31883 <= LPM_d0_ivl_31887(0 + 1 downto 0);
  tmp_ivl_31888 <= new_AGEMA_signal_3828 & n4098;
  LPM_q_ivl_31891 <= tmp_ivl_31893 & tmp_ivl_31888;
  tmp_ivl_31895 <= new_AGEMA_signal_3829 & n4210;
  LPM_q_ivl_31898 <= tmp_ivl_31900 & tmp_ivl_31895;
  tmp_ivl_31902 <= tmp_ivl_31906(1);
  tmp_ivl_31904 <= tmp_ivl_31906(0);
  tmp_ivl_31906 <= LPM_d0_ivl_31910(0 + 1 downto 0);
  tmp_ivl_31911 <= new_AGEMA_signal_3506 & n4099;
  LPM_q_ivl_31914 <= tmp_ivl_31916 & tmp_ivl_31911;
  tmp_ivl_31918 <= new_AGEMA_signal_4143 & n4228;
  LPM_q_ivl_31921 <= tmp_ivl_31923 & tmp_ivl_31918;
  new_AGEMA_signal_4435 <= tmp_ivl_31925(1);
  n4100 <= tmp_ivl_31925(0);
  tmp_ivl_31925 <= LPM_d0_ivl_31929(0 + 1 downto 0);
  tmp_ivl_31930 <= new_AGEMA_signal_3512 & n4101;
  LPM_q_ivl_31933 <= tmp_ivl_31935 & tmp_ivl_31930;
  tmp_ivl_31937 <= new_AGEMA_signal_4435 & n4100;
  LPM_q_ivl_31940 <= tmp_ivl_31942 & tmp_ivl_31937;
  new_AGEMA_signal_4566 <= tmp_ivl_31944(1);
  n4102 <= tmp_ivl_31944(0);
  tmp_ivl_31944 <= LPM_d0_ivl_31948(0 + 1 downto 0);
  tmp_ivl_31952 <= rcon(1);
  tmp_ivl_31953 <= tmp_ivl_31949 & tmp_ivl_31952;
  LPM_q_ivl_31956 <= tmp_ivl_31958 & tmp_ivl_31953;
  tmp_ivl_31960 <= new_AGEMA_signal_4566 & n4102;
  LPM_q_ivl_31963 <= tmp_ivl_31965 & tmp_ivl_31960;
  tmp_ivl_31967 <= tmp_ivl_31971(1);
  tmp_ivl_31969 <= tmp_ivl_31971(0);
  tmp_ivl_31971 <= LPM_d0_ivl_31975(0 + 1 downto 0);
  tmp_ivl_31976 <= new_AGEMA_signal_3502 & n4112;
  LPM_q_ivl_31979 <= tmp_ivl_31981 & tmp_ivl_31976;
  tmp_ivl_31983 <= new_AGEMA_signal_3511 & n4104;
  LPM_q_ivl_31986 <= tmp_ivl_31988 & tmp_ivl_31983;
  new_AGEMA_signal_3830 <= tmp_ivl_31990(1);
  n4105 <= tmp_ivl_31990(0);
  tmp_ivl_31990 <= LPM_d0_ivl_31994(0 + 1 downto 0);
  tmp_ivl_31995 <= new_AGEMA_signal_3503 & n4226;
  LPM_q_ivl_31998 <= tmp_ivl_32000 & tmp_ivl_31995;
  tmp_ivl_32002 <= new_AGEMA_signal_3830 & n4105;
  LPM_q_ivl_32005 <= tmp_ivl_32007 & tmp_ivl_32002;
  tmp_ivl_32009 <= tmp_ivl_32013(1);
  tmp_ivl_32011 <= tmp_ivl_32013(0);
  tmp_ivl_32013 <= LPM_d0_ivl_32017(0 + 1 downto 0);
  tmp_ivl_32018 <= new_AGEMA_signal_3502 & n4112;
  LPM_q_ivl_32021 <= tmp_ivl_32023 & tmp_ivl_32018;
  tmp_ivl_32025 <= new_AGEMA_signal_3501 & n4114;
  LPM_q_ivl_32028 <= tmp_ivl_32030 & tmp_ivl_32025;
  new_AGEMA_signal_3831 <= tmp_ivl_32032(1);
  n4106 <= tmp_ivl_32032(0);
  tmp_ivl_32032 <= LPM_d0_ivl_32036(0 + 1 downto 0);
  tmp_ivl_32037 <= new_AGEMA_signal_3509 & n4107;
  LPM_q_ivl_32040 <= tmp_ivl_32042 & tmp_ivl_32037;
  tmp_ivl_32044 <= new_AGEMA_signal_3831 & n4106;
  LPM_q_ivl_32047 <= tmp_ivl_32049 & tmp_ivl_32044;
  tmp_ivl_32051 <= tmp_ivl_32055(1);
  tmp_ivl_32053 <= tmp_ivl_32055(0);
  tmp_ivl_32055 <= LPM_d0_ivl_32059(0 + 1 downto 0);
  tmp_ivl_32060 <= new_AGEMA_signal_3508 & n4215;
  LPM_q_ivl_32063 <= tmp_ivl_32065 & tmp_ivl_32060;
  tmp_ivl_32067 <= new_AGEMA_signal_3501 & n4114;
  LPM_q_ivl_32070 <= tmp_ivl_32072 & tmp_ivl_32067;
  new_AGEMA_signal_3832 <= tmp_ivl_32074(1);
  n4108 <= tmp_ivl_32074(0);
  tmp_ivl_32074 <= LPM_d0_ivl_32078(0 + 1 downto 0);
  tmp_ivl_32079 <= new_AGEMA_signal_3500 & n4117;
  LPM_q_ivl_32082 <= tmp_ivl_32084 & tmp_ivl_32079;
  tmp_ivl_32086 <= new_AGEMA_signal_3832 & n4108;
  LPM_q_ivl_32089 <= tmp_ivl_32091 & tmp_ivl_32086;
  tmp_ivl_32093 <= tmp_ivl_32097(1);
  tmp_ivl_32095 <= tmp_ivl_32097(0);
  tmp_ivl_32097 <= LPM_d0_ivl_32101(0 + 1 downto 0);
  tmp_ivl_32102 <= new_AGEMA_signal_3499 & n4118;
  LPM_q_ivl_32105 <= tmp_ivl_32107 & tmp_ivl_32102;
  tmp_ivl_32109 <= new_AGEMA_signal_3505 & n4220;
  LPM_q_ivl_32112 <= tmp_ivl_32114 & tmp_ivl_32109;
  new_AGEMA_signal_3833 <= tmp_ivl_32116(1);
  n4109 <= tmp_ivl_32116(0);
  tmp_ivl_32116 <= LPM_d0_ivl_32120(0 + 1 downto 0);
  tmp_ivl_32121 <= new_AGEMA_signal_3500 & n4117;
  LPM_q_ivl_32124 <= tmp_ivl_32126 & tmp_ivl_32121;
  tmp_ivl_32128 <= new_AGEMA_signal_3833 & n4109;
  LPM_q_ivl_32131 <= tmp_ivl_32133 & tmp_ivl_32128;
  tmp_ivl_32135 <= tmp_ivl_32139(1);
  tmp_ivl_32137 <= tmp_ivl_32139(0);
  tmp_ivl_32139 <= LPM_d0_ivl_32143(0 + 1 downto 0);
  tmp_ivl_32144 <= new_AGEMA_signal_3499 & n4118;
  LPM_q_ivl_32147 <= tmp_ivl_32149 & tmp_ivl_32144;
  tmp_ivl_32151 <= new_AGEMA_signal_3504 & n4223;
  LPM_q_ivl_32154 <= tmp_ivl_32156 & tmp_ivl_32151;
  new_AGEMA_signal_3834 <= tmp_ivl_32158(1);
  n4110 <= tmp_ivl_32158(0);
  tmp_ivl_32158 <= LPM_d0_ivl_32162(0 + 1 downto 0);
  tmp_ivl_32163 <= new_AGEMA_signal_3498 & n4120;
  LPM_q_ivl_32166 <= tmp_ivl_32168 & tmp_ivl_32163;
  tmp_ivl_32170 <= new_AGEMA_signal_3834 & n4110;
  LPM_q_ivl_32173 <= tmp_ivl_32175 & tmp_ivl_32170;
  tmp_ivl_32177 <= tmp_ivl_32181(1);
  tmp_ivl_32179 <= tmp_ivl_32181(0);
  tmp_ivl_32181 <= LPM_d0_ivl_32185(0 + 1 downto 0);
  tmp_ivl_32186 <= new_AGEMA_signal_3498 & n4120;
  LPM_q_ivl_32189 <= tmp_ivl_32191 & tmp_ivl_32186;
  tmp_ivl_32193 <= new_AGEMA_signal_3497 & n4123;
  LPM_q_ivl_32196 <= tmp_ivl_32198 & tmp_ivl_32193;
  new_AGEMA_signal_3835 <= tmp_ivl_32200(1);
  n4111 <= tmp_ivl_32200(0);
  tmp_ivl_32200 <= LPM_d0_ivl_32204(0 + 1 downto 0);
  tmp_ivl_32205 <= new_AGEMA_signal_3503 & n4226;
  LPM_q_ivl_32208 <= tmp_ivl_32210 & tmp_ivl_32205;
  tmp_ivl_32212 <= new_AGEMA_signal_3835 & n4111;
  LPM_q_ivl_32215 <= tmp_ivl_32217 & tmp_ivl_32212;
  tmp_ivl_32219 <= tmp_ivl_32223(1);
  tmp_ivl_32221 <= tmp_ivl_32223(0);
  tmp_ivl_32223 <= LPM_d0_ivl_32227(0 + 1 downto 0);
  tmp_ivl_32228 <= new_AGEMA_signal_3502 & n4112;
  LPM_q_ivl_32231 <= tmp_ivl_32233 & tmp_ivl_32228;
  tmp_ivl_32235 <= new_AGEMA_signal_3496 & n4125;
  LPM_q_ivl_32238 <= tmp_ivl_32240 & tmp_ivl_32235;
  new_AGEMA_signal_3836 <= tmp_ivl_32242(1);
  n4113 <= tmp_ivl_32242(0);
  tmp_ivl_32242 <= LPM_d0_ivl_32246(0 + 1 downto 0);
  tmp_ivl_32247 <= new_AGEMA_signal_3497 & n4123;
  LPM_q_ivl_32250 <= tmp_ivl_32252 & tmp_ivl_32247;
  tmp_ivl_32254 <= new_AGEMA_signal_3836 & n4113;
  LPM_q_ivl_32257 <= tmp_ivl_32259 & tmp_ivl_32254;
  tmp_ivl_32261 <= tmp_ivl_32265(1);
  tmp_ivl_32263 <= tmp_ivl_32265(0);
  tmp_ivl_32265 <= LPM_d0_ivl_32269(0 + 1 downto 0);
  tmp_ivl_32270 <= new_AGEMA_signal_3495 & n4126;
  LPM_q_ivl_32273 <= tmp_ivl_32275 & tmp_ivl_32270;
  tmp_ivl_32277 <= new_AGEMA_signal_3501 & n4114;
  LPM_q_ivl_32280 <= tmp_ivl_32282 & tmp_ivl_32277;
  new_AGEMA_signal_3837 <= tmp_ivl_32284(1);
  n4115 <= tmp_ivl_32284(0);
  tmp_ivl_32284 <= LPM_d0_ivl_32288(0 + 1 downto 0);
  tmp_ivl_32289 <= new_AGEMA_signal_3496 & n4125;
  LPM_q_ivl_32292 <= tmp_ivl_32294 & tmp_ivl_32289;
  tmp_ivl_32296 <= new_AGEMA_signal_3837 & n4115;
  LPM_q_ivl_32299 <= tmp_ivl_32301 & tmp_ivl_32296;
  tmp_ivl_32303 <= tmp_ivl_32307(1);
  tmp_ivl_32305 <= tmp_ivl_32307(0);
  tmp_ivl_32307 <= LPM_d0_ivl_32311(0 + 1 downto 0);
  tmp_ivl_32312 <= new_AGEMA_signal_3495 & n4126;
  LPM_q_ivl_32315 <= tmp_ivl_32317 & tmp_ivl_32312;
  tmp_ivl_32319 <= new_AGEMA_signal_3494 & n4128;
  LPM_q_ivl_32322 <= tmp_ivl_32324 & tmp_ivl_32319;
  new_AGEMA_signal_3838 <= tmp_ivl_32326(1);
  n4116 <= tmp_ivl_32326(0);
  tmp_ivl_32326 <= LPM_d0_ivl_32330(0 + 1 downto 0);
  tmp_ivl_32331 <= new_AGEMA_signal_3500 & n4117;
  LPM_q_ivl_32334 <= tmp_ivl_32336 & tmp_ivl_32331;
  tmp_ivl_32338 <= new_AGEMA_signal_3838 & n4116;
  LPM_q_ivl_32341 <= tmp_ivl_32343 & tmp_ivl_32338;
  tmp_ivl_32345 <= tmp_ivl_32349(1);
  tmp_ivl_32347 <= tmp_ivl_32349(0);
  tmp_ivl_32349 <= LPM_d0_ivl_32353(0 + 1 downto 0);
  tmp_ivl_32354 <= new_AGEMA_signal_3499 & n4118;
  LPM_q_ivl_32357 <= tmp_ivl_32359 & tmp_ivl_32354;
  tmp_ivl_32361 <= new_AGEMA_signal_3494 & n4128;
  LPM_q_ivl_32364 <= tmp_ivl_32366 & tmp_ivl_32361;
  new_AGEMA_signal_3839 <= tmp_ivl_32368(1);
  n4119 <= tmp_ivl_32368(0);
  tmp_ivl_32368 <= LPM_d0_ivl_32372(0 + 1 downto 0);
  tmp_ivl_32373 <= new_AGEMA_signal_3493 & n4131;
  LPM_q_ivl_32376 <= tmp_ivl_32378 & tmp_ivl_32373;
  tmp_ivl_32380 <= new_AGEMA_signal_3839 & n4119;
  LPM_q_ivl_32383 <= tmp_ivl_32385 & tmp_ivl_32380;
  tmp_ivl_32387 <= tmp_ivl_32391(1);
  tmp_ivl_32389 <= tmp_ivl_32391(0);
  tmp_ivl_32391 <= LPM_d0_ivl_32395(0 + 1 downto 0);
  tmp_ivl_32396 <= new_AGEMA_signal_3498 & n4120;
  LPM_q_ivl_32399 <= tmp_ivl_32401 & tmp_ivl_32396;
  tmp_ivl_32403 <= new_AGEMA_signal_3492 & n4133;
  LPM_q_ivl_32406 <= tmp_ivl_32408 & tmp_ivl_32403;
  new_AGEMA_signal_3840 <= tmp_ivl_32410(1);
  n4121 <= tmp_ivl_32410(0);
  tmp_ivl_32410 <= LPM_d0_ivl_32414(0 + 1 downto 0);
  tmp_ivl_32415 <= new_AGEMA_signal_3493 & n4131;
  LPM_q_ivl_32418 <= tmp_ivl_32420 & tmp_ivl_32415;
  tmp_ivl_32422 <= new_AGEMA_signal_3840 & n4121;
  LPM_q_ivl_32425 <= tmp_ivl_32427 & tmp_ivl_32422;
  tmp_ivl_32429 <= tmp_ivl_32433(1);
  tmp_ivl_32431 <= tmp_ivl_32433(0);
  tmp_ivl_32433 <= LPM_d0_ivl_32437(0 + 1 downto 0);
  tmp_ivl_32438 <= new_AGEMA_signal_3491 & n4135;
  LPM_q_ivl_32441 <= tmp_ivl_32443 & tmp_ivl_32438;
  tmp_ivl_32445 <= new_AGEMA_signal_3492 & n4133;
  LPM_q_ivl_32448 <= tmp_ivl_32450 & tmp_ivl_32445;
  new_AGEMA_signal_3841 <= tmp_ivl_32452(1);
  n4122 <= tmp_ivl_32452(0);
  tmp_ivl_32452 <= LPM_d0_ivl_32456(0 + 1 downto 0);
  tmp_ivl_32457 <= new_AGEMA_signal_3497 & n4123;
  LPM_q_ivl_32460 <= tmp_ivl_32462 & tmp_ivl_32457;
  tmp_ivl_32464 <= new_AGEMA_signal_3841 & n4122;
  LPM_q_ivl_32467 <= tmp_ivl_32469 & tmp_ivl_32464;
  tmp_ivl_32471 <= tmp_ivl_32475(1);
  tmp_ivl_32473 <= tmp_ivl_32475(0);
  tmp_ivl_32475 <= LPM_d0_ivl_32479(0 + 1 downto 0);
  tmp_ivl_32480 <= new_AGEMA_signal_3490 & n4137;
  LPM_q_ivl_32483 <= tmp_ivl_32485 & tmp_ivl_32480;
  tmp_ivl_32487 <= new_AGEMA_signal_3491 & n4135;
  LPM_q_ivl_32490 <= tmp_ivl_32492 & tmp_ivl_32487;
  new_AGEMA_signal_3842 <= tmp_ivl_32494(1);
  n4124 <= tmp_ivl_32494(0);
  tmp_ivl_32494 <= LPM_d0_ivl_32498(0 + 1 downto 0);
  tmp_ivl_32499 <= new_AGEMA_signal_3496 & n4125;
  LPM_q_ivl_32502 <= tmp_ivl_32504 & tmp_ivl_32499;
  tmp_ivl_32506 <= new_AGEMA_signal_3842 & n4124;
  LPM_q_ivl_32509 <= tmp_ivl_32511 & tmp_ivl_32506;
  tmp_ivl_32513 <= tmp_ivl_32517(1);
  tmp_ivl_32515 <= tmp_ivl_32517(0);
  tmp_ivl_32517 <= LPM_d0_ivl_32521(0 + 1 downto 0);
  tmp_ivl_32522 <= new_AGEMA_signal_3495 & n4126;
  LPM_q_ivl_32525 <= tmp_ivl_32527 & tmp_ivl_32522;
  tmp_ivl_32529 <= new_AGEMA_signal_3489 & n4139;
  LPM_q_ivl_32532 <= tmp_ivl_32534 & tmp_ivl_32529;
  new_AGEMA_signal_3843 <= tmp_ivl_32536(1);
  n4127 <= tmp_ivl_32536(0);
  tmp_ivl_32536 <= LPM_d0_ivl_32540(0 + 1 downto 0);
  tmp_ivl_32541 <= new_AGEMA_signal_3490 & n4137;
  LPM_q_ivl_32544 <= tmp_ivl_32546 & tmp_ivl_32541;
  tmp_ivl_32548 <= new_AGEMA_signal_3843 & n4127;
  LPM_q_ivl_32551 <= tmp_ivl_32553 & tmp_ivl_32548;
  tmp_ivl_32555 <= tmp_ivl_32559(1);
  tmp_ivl_32557 <= tmp_ivl_32559(0);
  tmp_ivl_32559 <= LPM_d0_ivl_32563(0 + 1 downto 0);
  tmp_ivl_32564 <= new_AGEMA_signal_3494 & n4128;
  LPM_q_ivl_32567 <= tmp_ivl_32569 & tmp_ivl_32564;
  tmp_ivl_32571 <= new_AGEMA_signal_3488 & n4141;
  LPM_q_ivl_32574 <= tmp_ivl_32576 & tmp_ivl_32571;
  new_AGEMA_signal_3844 <= tmp_ivl_32578(1);
  n4129 <= tmp_ivl_32578(0);
  tmp_ivl_32578 <= LPM_d0_ivl_32582(0 + 1 downto 0);
  tmp_ivl_32583 <= new_AGEMA_signal_3489 & n4139;
  LPM_q_ivl_32586 <= tmp_ivl_32588 & tmp_ivl_32583;
  tmp_ivl_32590 <= new_AGEMA_signal_3844 & n4129;
  LPM_q_ivl_32593 <= tmp_ivl_32595 & tmp_ivl_32590;
  tmp_ivl_32597 <= tmp_ivl_32601(1);
  tmp_ivl_32599 <= tmp_ivl_32601(0);
  tmp_ivl_32601 <= LPM_d0_ivl_32605(0 + 1 downto 0);
  tmp_ivl_32606 <= new_AGEMA_signal_3487 & n4143;
  LPM_q_ivl_32609 <= tmp_ivl_32611 & tmp_ivl_32606;
  tmp_ivl_32613 <= new_AGEMA_signal_3488 & n4141;
  LPM_q_ivl_32616 <= tmp_ivl_32618 & tmp_ivl_32613;
  new_AGEMA_signal_3845 <= tmp_ivl_32620(1);
  n4130 <= tmp_ivl_32620(0);
  tmp_ivl_32620 <= LPM_d0_ivl_32624(0 + 1 downto 0);
  tmp_ivl_32625 <= new_AGEMA_signal_3493 & n4131;
  LPM_q_ivl_32628 <= tmp_ivl_32630 & tmp_ivl_32625;
  tmp_ivl_32632 <= new_AGEMA_signal_3845 & n4130;
  LPM_q_ivl_32635 <= tmp_ivl_32637 & tmp_ivl_32632;
  tmp_ivl_32639 <= tmp_ivl_32643(1);
  tmp_ivl_32641 <= tmp_ivl_32643(0);
  tmp_ivl_32643 <= LPM_d0_ivl_32647(0 + 1 downto 0);
  tmp_ivl_32648 <= new_AGEMA_signal_3486 & n4145;
  LPM_q_ivl_32651 <= tmp_ivl_32653 & tmp_ivl_32648;
  tmp_ivl_32655 <= new_AGEMA_signal_3487 & n4143;
  LPM_q_ivl_32658 <= tmp_ivl_32660 & tmp_ivl_32655;
  new_AGEMA_signal_3846 <= tmp_ivl_32662(1);
  n4132 <= tmp_ivl_32662(0);
  tmp_ivl_32662 <= LPM_d0_ivl_32666(0 + 1 downto 0);
  tmp_ivl_32667 <= new_AGEMA_signal_3492 & n4133;
  LPM_q_ivl_32670 <= tmp_ivl_32672 & tmp_ivl_32667;
  tmp_ivl_32674 <= new_AGEMA_signal_3846 & n4132;
  LPM_q_ivl_32677 <= tmp_ivl_32679 & tmp_ivl_32674;
  tmp_ivl_32681 <= tmp_ivl_32685(1);
  tmp_ivl_32683 <= tmp_ivl_32685(0);
  tmp_ivl_32685 <= LPM_d0_ivl_32689(0 + 1 downto 0);
  tmp_ivl_32690 <= new_AGEMA_signal_3485 & n4147;
  LPM_q_ivl_32693 <= tmp_ivl_32695 & tmp_ivl_32690;
  tmp_ivl_32697 <= new_AGEMA_signal_3486 & n4145;
  LPM_q_ivl_32700 <= tmp_ivl_32702 & tmp_ivl_32697;
  new_AGEMA_signal_3847 <= tmp_ivl_32704(1);
  n4134 <= tmp_ivl_32704(0);
  tmp_ivl_32704 <= LPM_d0_ivl_32708(0 + 1 downto 0);
  tmp_ivl_32709 <= new_AGEMA_signal_3491 & n4135;
  LPM_q_ivl_32712 <= tmp_ivl_32714 & tmp_ivl_32709;
  tmp_ivl_32716 <= new_AGEMA_signal_3847 & n4134;
  LPM_q_ivl_32719 <= tmp_ivl_32721 & tmp_ivl_32716;
  tmp_ivl_32723 <= tmp_ivl_32727(1);
  tmp_ivl_32725 <= tmp_ivl_32727(0);
  tmp_ivl_32727 <= LPM_d0_ivl_32731(0 + 1 downto 0);
  tmp_ivl_32732 <= new_AGEMA_signal_3484 & n4149;
  LPM_q_ivl_32735 <= tmp_ivl_32737 & tmp_ivl_32732;
  tmp_ivl_32739 <= new_AGEMA_signal_3485 & n4147;
  LPM_q_ivl_32742 <= tmp_ivl_32744 & tmp_ivl_32739;
  new_AGEMA_signal_3848 <= tmp_ivl_32746(1);
  n4136 <= tmp_ivl_32746(0);
  tmp_ivl_32746 <= LPM_d0_ivl_32750(0 + 1 downto 0);
  tmp_ivl_32751 <= new_AGEMA_signal_3490 & n4137;
  LPM_q_ivl_32754 <= tmp_ivl_32756 & tmp_ivl_32751;
  tmp_ivl_32758 <= new_AGEMA_signal_3848 & n4136;
  LPM_q_ivl_32761 <= tmp_ivl_32763 & tmp_ivl_32758;
  tmp_ivl_32765 <= tmp_ivl_32769(1);
  tmp_ivl_32767 <= tmp_ivl_32769(0);
  tmp_ivl_32769 <= LPM_d0_ivl_32773(0 + 1 downto 0);
  tmp_ivl_32774 <= new_AGEMA_signal_3483 & n4151;
  LPM_q_ivl_32777 <= tmp_ivl_32779 & tmp_ivl_32774;
  tmp_ivl_32781 <= new_AGEMA_signal_3484 & n4149;
  LPM_q_ivl_32784 <= tmp_ivl_32786 & tmp_ivl_32781;
  new_AGEMA_signal_3849 <= tmp_ivl_32788(1);
  n4138 <= tmp_ivl_32788(0);
  tmp_ivl_32788 <= LPM_d0_ivl_32792(0 + 1 downto 0);
  tmp_ivl_32793 <= new_AGEMA_signal_3489 & n4139;
  LPM_q_ivl_32796 <= tmp_ivl_32798 & tmp_ivl_32793;
  tmp_ivl_32800 <= new_AGEMA_signal_3849 & n4138;
  LPM_q_ivl_32803 <= tmp_ivl_32805 & tmp_ivl_32800;
  tmp_ivl_32807 <= tmp_ivl_32811(1);
  tmp_ivl_32809 <= tmp_ivl_32811(0);
  tmp_ivl_32811 <= LPM_d0_ivl_32815(0 + 1 downto 0);
  tmp_ivl_32816 <= new_AGEMA_signal_3482 & n4153;
  LPM_q_ivl_32819 <= tmp_ivl_32821 & tmp_ivl_32816;
  tmp_ivl_32823 <= new_AGEMA_signal_3483 & n4151;
  LPM_q_ivl_32826 <= tmp_ivl_32828 & tmp_ivl_32823;
  new_AGEMA_signal_3850 <= tmp_ivl_32830(1);
  n4140 <= tmp_ivl_32830(0);
  tmp_ivl_32830 <= LPM_d0_ivl_32834(0 + 1 downto 0);
  tmp_ivl_32835 <= new_AGEMA_signal_3488 & n4141;
  LPM_q_ivl_32838 <= tmp_ivl_32840 & tmp_ivl_32835;
  tmp_ivl_32842 <= new_AGEMA_signal_3850 & n4140;
  LPM_q_ivl_32845 <= tmp_ivl_32847 & tmp_ivl_32842;
  tmp_ivl_32849 <= tmp_ivl_32853(1);
  tmp_ivl_32851 <= tmp_ivl_32853(0);
  tmp_ivl_32853 <= LPM_d0_ivl_32857(0 + 1 downto 0);
  tmp_ivl_32858 <= new_AGEMA_signal_3481 & n4155;
  LPM_q_ivl_32861 <= tmp_ivl_32863 & tmp_ivl_32858;
  tmp_ivl_32865 <= new_AGEMA_signal_3482 & n4153;
  LPM_q_ivl_32868 <= tmp_ivl_32870 & tmp_ivl_32865;
  new_AGEMA_signal_3851 <= tmp_ivl_32872(1);
  n4142 <= tmp_ivl_32872(0);
  tmp_ivl_32872 <= LPM_d0_ivl_32876(0 + 1 downto 0);
  tmp_ivl_32877 <= new_AGEMA_signal_3487 & n4143;
  LPM_q_ivl_32880 <= tmp_ivl_32882 & tmp_ivl_32877;
  tmp_ivl_32884 <= new_AGEMA_signal_3851 & n4142;
  LPM_q_ivl_32887 <= tmp_ivl_32889 & tmp_ivl_32884;
  tmp_ivl_32891 <= tmp_ivl_32895(1);
  tmp_ivl_32893 <= tmp_ivl_32895(0);
  tmp_ivl_32895 <= LPM_d0_ivl_32899(0 + 1 downto 0);
  tmp_ivl_32900 <= new_AGEMA_signal_3480 & n4157;
  LPM_q_ivl_32903 <= tmp_ivl_32905 & tmp_ivl_32900;
  tmp_ivl_32907 <= new_AGEMA_signal_3481 & n4155;
  LPM_q_ivl_32910 <= tmp_ivl_32912 & tmp_ivl_32907;
  new_AGEMA_signal_3852 <= tmp_ivl_32914(1);
  n4144 <= tmp_ivl_32914(0);
  tmp_ivl_32914 <= LPM_d0_ivl_32918(0 + 1 downto 0);
  tmp_ivl_32919 <= new_AGEMA_signal_3486 & n4145;
  LPM_q_ivl_32922 <= tmp_ivl_32924 & tmp_ivl_32919;
  tmp_ivl_32926 <= new_AGEMA_signal_3852 & n4144;
  LPM_q_ivl_32929 <= tmp_ivl_32931 & tmp_ivl_32926;
  tmp_ivl_32933 <= tmp_ivl_32937(1);
  tmp_ivl_32935 <= tmp_ivl_32937(0);
  tmp_ivl_32937 <= LPM_d0_ivl_32941(0 + 1 downto 0);
  tmp_ivl_32942 <= new_AGEMA_signal_3478 & n4159;
  LPM_q_ivl_32945 <= tmp_ivl_32947 & tmp_ivl_32942;
  tmp_ivl_32949 <= new_AGEMA_signal_3480 & n4157;
  LPM_q_ivl_32952 <= tmp_ivl_32954 & tmp_ivl_32949;
  new_AGEMA_signal_3853 <= tmp_ivl_32956(1);
  n4146 <= tmp_ivl_32956(0);
  tmp_ivl_32956 <= LPM_d0_ivl_32960(0 + 1 downto 0);
  tmp_ivl_32961 <= new_AGEMA_signal_3485 & n4147;
  LPM_q_ivl_32964 <= tmp_ivl_32966 & tmp_ivl_32961;
  tmp_ivl_32968 <= new_AGEMA_signal_3853 & n4146;
  LPM_q_ivl_32971 <= tmp_ivl_32973 & tmp_ivl_32968;
  tmp_ivl_32975 <= tmp_ivl_32979(1);
  tmp_ivl_32977 <= tmp_ivl_32979(0);
  tmp_ivl_32979 <= LPM_d0_ivl_32983(0 + 1 downto 0);
  tmp_ivl_32984 <= new_AGEMA_signal_3476 & n4161;
  LPM_q_ivl_32987 <= tmp_ivl_32989 & tmp_ivl_32984;
  tmp_ivl_32991 <= new_AGEMA_signal_3478 & n4159;
  LPM_q_ivl_32994 <= tmp_ivl_32996 & tmp_ivl_32991;
  new_AGEMA_signal_3854 <= tmp_ivl_32998(1);
  n4148 <= tmp_ivl_32998(0);
  tmp_ivl_32998 <= LPM_d0_ivl_33002(0 + 1 downto 0);
  tmp_ivl_33003 <= new_AGEMA_signal_3484 & n4149;
  LPM_q_ivl_33006 <= tmp_ivl_33008 & tmp_ivl_33003;
  tmp_ivl_33010 <= new_AGEMA_signal_3854 & n4148;
  LPM_q_ivl_33013 <= tmp_ivl_33015 & tmp_ivl_33010;
  tmp_ivl_33017 <= tmp_ivl_33021(1);
  tmp_ivl_33019 <= tmp_ivl_33021(0);
  tmp_ivl_33021 <= LPM_d0_ivl_33025(0 + 1 downto 0);
  tmp_ivl_33026 <= new_AGEMA_signal_3474 & n4163;
  LPM_q_ivl_33029 <= tmp_ivl_33031 & tmp_ivl_33026;
  tmp_ivl_33033 <= new_AGEMA_signal_3476 & n4161;
  LPM_q_ivl_33036 <= tmp_ivl_33038 & tmp_ivl_33033;
  new_AGEMA_signal_3855 <= tmp_ivl_33040(1);
  n4150 <= tmp_ivl_33040(0);
  tmp_ivl_33040 <= LPM_d0_ivl_33044(0 + 1 downto 0);
  tmp_ivl_33045 <= new_AGEMA_signal_3483 & n4151;
  LPM_q_ivl_33048 <= tmp_ivl_33050 & tmp_ivl_33045;
  tmp_ivl_33052 <= new_AGEMA_signal_3855 & n4150;
  LPM_q_ivl_33055 <= tmp_ivl_33057 & tmp_ivl_33052;
  tmp_ivl_33059 <= tmp_ivl_33063(1);
  tmp_ivl_33061 <= tmp_ivl_33063(0);
  tmp_ivl_33063 <= LPM_d0_ivl_33067(0 + 1 downto 0);
  tmp_ivl_33068 <= new_AGEMA_signal_3471 & n4164;
  LPM_q_ivl_33071 <= tmp_ivl_33073 & tmp_ivl_33068;
  tmp_ivl_33075 <= new_AGEMA_signal_3474 & n4163;
  LPM_q_ivl_33078 <= tmp_ivl_33080 & tmp_ivl_33075;
  new_AGEMA_signal_3856 <= tmp_ivl_33082(1);
  n4152 <= tmp_ivl_33082(0);
  tmp_ivl_33082 <= LPM_d0_ivl_33086(0 + 1 downto 0);
  tmp_ivl_33087 <= new_AGEMA_signal_3482 & n4153;
  LPM_q_ivl_33090 <= tmp_ivl_33092 & tmp_ivl_33087;
  tmp_ivl_33094 <= new_AGEMA_signal_3856 & n4152;
  LPM_q_ivl_33097 <= tmp_ivl_33099 & tmp_ivl_33094;
  tmp_ivl_33101 <= tmp_ivl_33105(1);
  tmp_ivl_33103 <= tmp_ivl_33105(0);
  tmp_ivl_33105 <= LPM_d0_ivl_33109(0 + 1 downto 0);
  tmp_ivl_33110 <= new_AGEMA_signal_3468 & n4166;
  LPM_q_ivl_33113 <= tmp_ivl_33115 & tmp_ivl_33110;
  tmp_ivl_33117 <= new_AGEMA_signal_3471 & n4164;
  LPM_q_ivl_33120 <= tmp_ivl_33122 & tmp_ivl_33117;
  new_AGEMA_signal_3857 <= tmp_ivl_33124(1);
  n4154 <= tmp_ivl_33124(0);
  tmp_ivl_33124 <= LPM_d0_ivl_33128(0 + 1 downto 0);
  tmp_ivl_33129 <= new_AGEMA_signal_3481 & n4155;
  LPM_q_ivl_33132 <= tmp_ivl_33134 & tmp_ivl_33129;
  tmp_ivl_33136 <= new_AGEMA_signal_3857 & n4154;
  LPM_q_ivl_33139 <= tmp_ivl_33141 & tmp_ivl_33136;
  tmp_ivl_33143 <= tmp_ivl_33147(1);
  tmp_ivl_33145 <= tmp_ivl_33147(0);
  tmp_ivl_33147 <= LPM_d0_ivl_33151(0 + 1 downto 0);
  tmp_ivl_33152 <= new_AGEMA_signal_3465 & n4169;
  LPM_q_ivl_33155 <= tmp_ivl_33157 & tmp_ivl_33152;
  tmp_ivl_33159 <= new_AGEMA_signal_3468 & n4166;
  LPM_q_ivl_33162 <= tmp_ivl_33164 & tmp_ivl_33159;
  new_AGEMA_signal_3858 <= tmp_ivl_33166(1);
  n4156 <= tmp_ivl_33166(0);
  tmp_ivl_33166 <= LPM_d0_ivl_33170(0 + 1 downto 0);
  tmp_ivl_33171 <= new_AGEMA_signal_3480 & n4157;
  LPM_q_ivl_33174 <= tmp_ivl_33176 & tmp_ivl_33171;
  tmp_ivl_33178 <= new_AGEMA_signal_3858 & n4156;
  LPM_q_ivl_33181 <= tmp_ivl_33183 & tmp_ivl_33178;
  tmp_ivl_33185 <= tmp_ivl_33189(1);
  tmp_ivl_33187 <= tmp_ivl_33189(0);
  tmp_ivl_33189 <= LPM_d0_ivl_33193(0 + 1 downto 0);
  tmp_ivl_33194 <= new_AGEMA_signal_3462 & n4170;
  LPM_q_ivl_33197 <= tmp_ivl_33199 & tmp_ivl_33194;
  tmp_ivl_33201 <= new_AGEMA_signal_3465 & n4169;
  LPM_q_ivl_33204 <= tmp_ivl_33206 & tmp_ivl_33201;
  new_AGEMA_signal_3859 <= tmp_ivl_33208(1);
  n4158 <= tmp_ivl_33208(0);
  tmp_ivl_33208 <= LPM_d0_ivl_33212(0 + 1 downto 0);
  tmp_ivl_33213 <= new_AGEMA_signal_3478 & n4159;
  LPM_q_ivl_33216 <= tmp_ivl_33218 & tmp_ivl_33213;
  tmp_ivl_33220 <= new_AGEMA_signal_3859 & n4158;
  LPM_q_ivl_33223 <= tmp_ivl_33225 & tmp_ivl_33220;
  tmp_ivl_33227 <= tmp_ivl_33231(1);
  tmp_ivl_33229 <= tmp_ivl_33231(0);
  tmp_ivl_33231 <= LPM_d0_ivl_33235(0 + 1 downto 0);
  tmp_ivl_33236 <= new_AGEMA_signal_3459 & n4172;
  LPM_q_ivl_33239 <= tmp_ivl_33241 & tmp_ivl_33236;
  tmp_ivl_33243 <= new_AGEMA_signal_3462 & n4170;
  LPM_q_ivl_33246 <= tmp_ivl_33248 & tmp_ivl_33243;
  new_AGEMA_signal_3860 <= tmp_ivl_33250(1);
  n4160 <= tmp_ivl_33250(0);
  tmp_ivl_33250 <= LPM_d0_ivl_33254(0 + 1 downto 0);
  tmp_ivl_33255 <= new_AGEMA_signal_3476 & n4161;
  LPM_q_ivl_33258 <= tmp_ivl_33260 & tmp_ivl_33255;
  tmp_ivl_33262 <= new_AGEMA_signal_3860 & n4160;
  LPM_q_ivl_33265 <= tmp_ivl_33267 & tmp_ivl_33262;
  tmp_ivl_33269 <= tmp_ivl_33273(1);
  tmp_ivl_33271 <= tmp_ivl_33273(0);
  tmp_ivl_33273 <= LPM_d0_ivl_33277(0 + 1 downto 0);
  tmp_ivl_33278 <= new_AGEMA_signal_3456 & n4174;
  LPM_q_ivl_33281 <= tmp_ivl_33283 & tmp_ivl_33278;
  tmp_ivl_33285 <= new_AGEMA_signal_3459 & n4172;
  LPM_q_ivl_33288 <= tmp_ivl_33290 & tmp_ivl_33285;
  new_AGEMA_signal_3861 <= tmp_ivl_33292(1);
  n4162 <= tmp_ivl_33292(0);
  tmp_ivl_33292 <= LPM_d0_ivl_33296(0 + 1 downto 0);
  tmp_ivl_33297 <= new_AGEMA_signal_3474 & n4163;
  LPM_q_ivl_33300 <= tmp_ivl_33302 & tmp_ivl_33297;
  tmp_ivl_33304 <= new_AGEMA_signal_3861 & n4162;
  LPM_q_ivl_33307 <= tmp_ivl_33309 & tmp_ivl_33304;
  tmp_ivl_33311 <= tmp_ivl_33315(1);
  tmp_ivl_33313 <= tmp_ivl_33315(0);
  tmp_ivl_33315 <= LPM_d0_ivl_33319(0 + 1 downto 0);
  tmp_ivl_33320 <= new_AGEMA_signal_3456 & n4174;
  LPM_q_ivl_33323 <= tmp_ivl_33325 & tmp_ivl_33320;
  tmp_ivl_33327 <= new_AGEMA_signal_3471 & n4164;
  LPM_q_ivl_33330 <= tmp_ivl_33332 & tmp_ivl_33327;
  new_AGEMA_signal_3862 <= tmp_ivl_33334(1);
  n4165 <= tmp_ivl_33334(0);
  tmp_ivl_33334 <= LPM_d0_ivl_33338(0 + 1 downto 0);
  tmp_ivl_33339 <= new_AGEMA_signal_3473 & n4177;
  LPM_q_ivl_33342 <= tmp_ivl_33344 & tmp_ivl_33339;
  tmp_ivl_33346 <= new_AGEMA_signal_3862 & n4165;
  LPM_q_ivl_33349 <= tmp_ivl_33351 & tmp_ivl_33346;
  tmp_ivl_33353 <= tmp_ivl_33357(1);
  tmp_ivl_33355 <= tmp_ivl_33357(0);
  tmp_ivl_33357 <= LPM_d0_ivl_33361(0 + 1 downto 0);
  tmp_ivl_33362 <= new_AGEMA_signal_3470 & n4178;
  LPM_q_ivl_33365 <= tmp_ivl_33367 & tmp_ivl_33362;
  tmp_ivl_33369 <= new_AGEMA_signal_3468 & n4166;
  LPM_q_ivl_33372 <= tmp_ivl_33374 & tmp_ivl_33369;
  new_AGEMA_signal_3863 <= tmp_ivl_33376(1);
  n4167 <= tmp_ivl_33376(0);
  tmp_ivl_33376 <= LPM_d0_ivl_33380(0 + 1 downto 0);
  tmp_ivl_33381 <= new_AGEMA_signal_3473 & n4177;
  LPM_q_ivl_33384 <= tmp_ivl_33386 & tmp_ivl_33381;
  tmp_ivl_33388 <= new_AGEMA_signal_3863 & n4167;
  LPM_q_ivl_33391 <= tmp_ivl_33393 & tmp_ivl_33388;
  tmp_ivl_33395 <= tmp_ivl_33399(1);
  tmp_ivl_33397 <= tmp_ivl_33399(0);
  tmp_ivl_33399 <= LPM_d0_ivl_33403(0 + 1 downto 0);
  tmp_ivl_33404 <= new_AGEMA_signal_3470 & n4178;
  LPM_q_ivl_33407 <= tmp_ivl_33409 & tmp_ivl_33404;
  tmp_ivl_33411 <= new_AGEMA_signal_3466 & n4180;
  LPM_q_ivl_33414 <= tmp_ivl_33416 & tmp_ivl_33411;
  new_AGEMA_signal_3864 <= tmp_ivl_33418(1);
  n4168 <= tmp_ivl_33418(0);
  tmp_ivl_33418 <= LPM_d0_ivl_33422(0 + 1 downto 0);
  tmp_ivl_33423 <= new_AGEMA_signal_3465 & n4169;
  LPM_q_ivl_33426 <= tmp_ivl_33428 & tmp_ivl_33423;
  tmp_ivl_33430 <= new_AGEMA_signal_3864 & n4168;
  LPM_q_ivl_33433 <= tmp_ivl_33435 & tmp_ivl_33430;
  tmp_ivl_33437 <= tmp_ivl_33441(1);
  tmp_ivl_33439 <= tmp_ivl_33441(0);
  tmp_ivl_33441 <= LPM_d0_ivl_33445(0 + 1 downto 0);
  tmp_ivl_33446 <= new_AGEMA_signal_3466 & n4180;
  LPM_q_ivl_33449 <= tmp_ivl_33451 & tmp_ivl_33446;
  tmp_ivl_33453 <= new_AGEMA_signal_3462 & n4170;
  LPM_q_ivl_33456 <= tmp_ivl_33458 & tmp_ivl_33453;
  new_AGEMA_signal_3865 <= tmp_ivl_33460(1);
  n4171 <= tmp_ivl_33460(0);
  tmp_ivl_33460 <= LPM_d0_ivl_33464(0 + 1 downto 0);
  tmp_ivl_33465 <= new_AGEMA_signal_3464 & n4183;
  LPM_q_ivl_33468 <= tmp_ivl_33470 & tmp_ivl_33465;
  tmp_ivl_33472 <= new_AGEMA_signal_3865 & n4171;
  LPM_q_ivl_33475 <= tmp_ivl_33477 & tmp_ivl_33472;
  tmp_ivl_33479 <= tmp_ivl_33483(1);
  tmp_ivl_33481 <= tmp_ivl_33483(0);
  tmp_ivl_33483 <= LPM_d0_ivl_33487(0 + 1 downto 0);
  tmp_ivl_33488 <= new_AGEMA_signal_3459 & n4172;
  LPM_q_ivl_33491 <= tmp_ivl_33493 & tmp_ivl_33488;
  tmp_ivl_33495 <= new_AGEMA_signal_3461 & n4184;
  LPM_q_ivl_33498 <= tmp_ivl_33500 & tmp_ivl_33495;
  new_AGEMA_signal_3866 <= tmp_ivl_33502(1);
  n4173 <= tmp_ivl_33502(0);
  tmp_ivl_33502 <= LPM_d0_ivl_33506(0 + 1 downto 0);
  tmp_ivl_33507 <= new_AGEMA_signal_3464 & n4183;
  LPM_q_ivl_33510 <= tmp_ivl_33512 & tmp_ivl_33507;
  tmp_ivl_33514 <= new_AGEMA_signal_3866 & n4173;
  LPM_q_ivl_33517 <= tmp_ivl_33519 & tmp_ivl_33514;
  tmp_ivl_33521 <= tmp_ivl_33525(1);
  tmp_ivl_33523 <= tmp_ivl_33525(0);
  tmp_ivl_33525 <= LPM_d0_ivl_33529(0 + 1 downto 0);
  tmp_ivl_33530 <= new_AGEMA_signal_3457 & n4186;
  LPM_q_ivl_33533 <= tmp_ivl_33535 & tmp_ivl_33530;
  tmp_ivl_33537 <= new_AGEMA_signal_3456 & n4174;
  LPM_q_ivl_33540 <= tmp_ivl_33542 & tmp_ivl_33537;
  new_AGEMA_signal_3867 <= tmp_ivl_33544(1);
  n4175 <= tmp_ivl_33544(0);
  tmp_ivl_33544 <= LPM_d0_ivl_33548(0 + 1 downto 0);
  tmp_ivl_33549 <= new_AGEMA_signal_3461 & n4184;
  LPM_q_ivl_33552 <= tmp_ivl_33554 & tmp_ivl_33549;
  tmp_ivl_33556 <= new_AGEMA_signal_3867 & n4175;
  LPM_q_ivl_33559 <= tmp_ivl_33561 & tmp_ivl_33556;
  tmp_ivl_33563 <= tmp_ivl_33567(1);
  tmp_ivl_33565 <= tmp_ivl_33567(0);
  tmp_ivl_33567 <= LPM_d0_ivl_33571(0 + 1 downto 0);
  tmp_ivl_33572 <= new_AGEMA_signal_3457 & n4186;
  LPM_q_ivl_33575 <= tmp_ivl_33577 & tmp_ivl_33572;
  tmp_ivl_33579 <= new_AGEMA_signal_3455 & n4189;
  LPM_q_ivl_33582 <= tmp_ivl_33584 & tmp_ivl_33579;
  new_AGEMA_signal_3868 <= tmp_ivl_33586(1);
  n4176 <= tmp_ivl_33586(0);
  tmp_ivl_33586 <= LPM_d0_ivl_33590(0 + 1 downto 0);
  tmp_ivl_33591 <= new_AGEMA_signal_3473 & n4177;
  LPM_q_ivl_33594 <= tmp_ivl_33596 & tmp_ivl_33591;
  tmp_ivl_33598 <= new_AGEMA_signal_3868 & n4176;
  LPM_q_ivl_33601 <= tmp_ivl_33603 & tmp_ivl_33598;
  tmp_ivl_33605 <= tmp_ivl_33609(1);
  tmp_ivl_33607 <= tmp_ivl_33609(0);
  tmp_ivl_33609 <= LPM_d0_ivl_33613(0 + 1 downto 0);
  tmp_ivl_33614 <= new_AGEMA_signal_3470 & n4178;
  LPM_q_ivl_33617 <= tmp_ivl_33619 & tmp_ivl_33614;
  tmp_ivl_33621 <= new_AGEMA_signal_3455 & n4189;
  LPM_q_ivl_33624 <= tmp_ivl_33626 & tmp_ivl_33621;
  new_AGEMA_signal_3869 <= tmp_ivl_33628(1);
  n4179 <= tmp_ivl_33628(0);
  tmp_ivl_33628 <= LPM_d0_ivl_33632(0 + 1 downto 0);
  tmp_ivl_33633 <= new_AGEMA_signal_3479 & n4191;
  LPM_q_ivl_33636 <= tmp_ivl_33638 & tmp_ivl_33633;
  tmp_ivl_33640 <= new_AGEMA_signal_3869 & n4179;
  LPM_q_ivl_33643 <= tmp_ivl_33645 & tmp_ivl_33640;
  tmp_ivl_33647 <= tmp_ivl_33651(1);
  tmp_ivl_33649 <= tmp_ivl_33651(0);
  tmp_ivl_33651 <= LPM_d0_ivl_33655(0 + 1 downto 0);
  tmp_ivl_33656 <= new_AGEMA_signal_3477 & n4193;
  LPM_q_ivl_33659 <= tmp_ivl_33661 & tmp_ivl_33656;
  tmp_ivl_33663 <= new_AGEMA_signal_3466 & n4180;
  LPM_q_ivl_33666 <= tmp_ivl_33668 & tmp_ivl_33663;
  new_AGEMA_signal_3870 <= tmp_ivl_33670(1);
  n4181 <= tmp_ivl_33670(0);
  tmp_ivl_33670 <= LPM_d0_ivl_33674(0 + 1 downto 0);
  tmp_ivl_33675 <= new_AGEMA_signal_3479 & n4191;
  LPM_q_ivl_33678 <= tmp_ivl_33680 & tmp_ivl_33675;
  tmp_ivl_33682 <= new_AGEMA_signal_3870 & n4181;
  LPM_q_ivl_33685 <= tmp_ivl_33687 & tmp_ivl_33682;
  tmp_ivl_33689 <= tmp_ivl_33693(1);
  tmp_ivl_33691 <= tmp_ivl_33693(0);
  tmp_ivl_33693 <= LPM_d0_ivl_33697(0 + 1 downto 0);
  tmp_ivl_33698 <= new_AGEMA_signal_3477 & n4193;
  LPM_q_ivl_33701 <= tmp_ivl_33703 & tmp_ivl_33698;
  tmp_ivl_33705 <= new_AGEMA_signal_3475 & n4195;
  LPM_q_ivl_33708 <= tmp_ivl_33710 & tmp_ivl_33705;
  new_AGEMA_signal_3871 <= tmp_ivl_33712(1);
  n4182 <= tmp_ivl_33712(0);
  tmp_ivl_33712 <= LPM_d0_ivl_33716(0 + 1 downto 0);
  tmp_ivl_33717 <= new_AGEMA_signal_3464 & n4183;
  LPM_q_ivl_33720 <= tmp_ivl_33722 & tmp_ivl_33717;
  tmp_ivl_33724 <= new_AGEMA_signal_3871 & n4182;
  LPM_q_ivl_33727 <= tmp_ivl_33729 & tmp_ivl_33724;
  tmp_ivl_33731 <= tmp_ivl_33735(1);
  tmp_ivl_33733 <= tmp_ivl_33735(0);
  tmp_ivl_33735 <= LPM_d0_ivl_33739(0 + 1 downto 0);
  tmp_ivl_33740 <= new_AGEMA_signal_3475 & n4195;
  LPM_q_ivl_33743 <= tmp_ivl_33745 & tmp_ivl_33740;
  tmp_ivl_33747 <= new_AGEMA_signal_3461 & n4184;
  LPM_q_ivl_33750 <= tmp_ivl_33752 & tmp_ivl_33747;
  new_AGEMA_signal_3872 <= tmp_ivl_33754(1);
  n4185 <= tmp_ivl_33754(0);
  tmp_ivl_33754 <= LPM_d0_ivl_33758(0 + 1 downto 0);
  tmp_ivl_33759 <= new_AGEMA_signal_3472 & n4198;
  LPM_q_ivl_33762 <= tmp_ivl_33764 & tmp_ivl_33759;
  tmp_ivl_33766 <= new_AGEMA_signal_3872 & n4185;
  LPM_q_ivl_33769 <= tmp_ivl_33771 & tmp_ivl_33766;
  tmp_ivl_33773 <= tmp_ivl_33777(1);
  tmp_ivl_33775 <= tmp_ivl_33777(0);
  tmp_ivl_33777 <= LPM_d0_ivl_33781(0 + 1 downto 0);
  tmp_ivl_33782 <= new_AGEMA_signal_3469 & n4199;
  LPM_q_ivl_33785 <= tmp_ivl_33787 & tmp_ivl_33782;
  tmp_ivl_33789 <= new_AGEMA_signal_3457 & n4186;
  LPM_q_ivl_33792 <= tmp_ivl_33794 & tmp_ivl_33789;
  new_AGEMA_signal_3873 <= tmp_ivl_33796(1);
  n4187 <= tmp_ivl_33796(0);
  tmp_ivl_33796 <= LPM_d0_ivl_33800(0 + 1 downto 0);
  tmp_ivl_33801 <= new_AGEMA_signal_3472 & n4198;
  LPM_q_ivl_33804 <= tmp_ivl_33806 & tmp_ivl_33801;
  tmp_ivl_33808 <= new_AGEMA_signal_3873 & n4187;
  LPM_q_ivl_33811 <= tmp_ivl_33813 & tmp_ivl_33808;
  tmp_ivl_33815 <= tmp_ivl_33819(1);
  tmp_ivl_33817 <= tmp_ivl_33819(0);
  tmp_ivl_33819 <= LPM_d0_ivl_33823(0 + 1 downto 0);
  tmp_ivl_33824 <= new_AGEMA_signal_3469 & n4199;
  LPM_q_ivl_33827 <= tmp_ivl_33829 & tmp_ivl_33824;
  tmp_ivl_33831 <= new_AGEMA_signal_3467 & n4201;
  LPM_q_ivl_33834 <= tmp_ivl_33836 & tmp_ivl_33831;
  new_AGEMA_signal_3874 <= tmp_ivl_33838(1);
  n4188 <= tmp_ivl_33838(0);
  tmp_ivl_33838 <= LPM_d0_ivl_33842(0 + 1 downto 0);
  tmp_ivl_33843 <= new_AGEMA_signal_3455 & n4189;
  LPM_q_ivl_33846 <= tmp_ivl_33848 & tmp_ivl_33843;
  tmp_ivl_33850 <= new_AGEMA_signal_3874 & n4188;
  LPM_q_ivl_33853 <= tmp_ivl_33855 & tmp_ivl_33850;
  tmp_ivl_33857 <= tmp_ivl_33861(1);
  tmp_ivl_33859 <= tmp_ivl_33861(0);
  tmp_ivl_33861 <= LPM_d0_ivl_33865(0 + 1 downto 0);
  tmp_ivl_33866 <= new_AGEMA_signal_3467 & n4201;
  LPM_q_ivl_33869 <= tmp_ivl_33871 & tmp_ivl_33866;
  tmp_ivl_33873 <= new_AGEMA_signal_3463 & n4192;
  LPM_q_ivl_33876 <= tmp_ivl_33878 & tmp_ivl_33873;
  new_AGEMA_signal_3875 <= tmp_ivl_33880(1);
  n4190 <= tmp_ivl_33880(0);
  tmp_ivl_33880 <= LPM_d0_ivl_33884(0 + 1 downto 0);
  tmp_ivl_33885 <= new_AGEMA_signal_3479 & n4191;
  LPM_q_ivl_33888 <= tmp_ivl_33890 & tmp_ivl_33885;
  tmp_ivl_33892 <= new_AGEMA_signal_3875 & n4190;
  LPM_q_ivl_33895 <= tmp_ivl_33897 & tmp_ivl_33892;
  tmp_ivl_33899 <= tmp_ivl_33903(1);
  tmp_ivl_33901 <= tmp_ivl_33903(0);
  tmp_ivl_33903 <= LPM_d0_ivl_33907(0 + 1 downto 0);
  tmp_ivl_33908 <= new_AGEMA_signal_3477 & n4193;
  LPM_q_ivl_33911 <= tmp_ivl_33913 & tmp_ivl_33908;
  tmp_ivl_33915 <= new_AGEMA_signal_3463 & n4192;
  LPM_q_ivl_33918 <= tmp_ivl_33920 & tmp_ivl_33915;
  new_AGEMA_signal_3876 <= tmp_ivl_33922(1);
  n4194 <= tmp_ivl_33922(0);
  tmp_ivl_33922 <= LPM_d0_ivl_33926(0 + 1 downto 0);
  tmp_ivl_33927 <= new_AGEMA_signal_3460 & n4204;
  LPM_q_ivl_33930 <= tmp_ivl_33932 & tmp_ivl_33927;
  tmp_ivl_33934 <= new_AGEMA_signal_3876 & n4194;
  LPM_q_ivl_33937 <= tmp_ivl_33939 & tmp_ivl_33934;
  tmp_ivl_33941 <= tmp_ivl_33945(1);
  tmp_ivl_33943 <= tmp_ivl_33945(0);
  tmp_ivl_33945 <= LPM_d0_ivl_33949(0 + 1 downto 0);
  tmp_ivl_33950 <= new_AGEMA_signal_3458 & n4212;
  LPM_q_ivl_33953 <= tmp_ivl_33955 & tmp_ivl_33950;
  tmp_ivl_33957 <= new_AGEMA_signal_3475 & n4195;
  LPM_q_ivl_33960 <= tmp_ivl_33962 & tmp_ivl_33957;
  new_AGEMA_signal_3877 <= tmp_ivl_33964(1);
  n4196 <= tmp_ivl_33964(0);
  tmp_ivl_33964 <= LPM_d0_ivl_33968(0 + 1 downto 0);
  tmp_ivl_33969 <= new_AGEMA_signal_3460 & n4204;
  LPM_q_ivl_33972 <= tmp_ivl_33974 & tmp_ivl_33969;
  tmp_ivl_33976 <= new_AGEMA_signal_3877 & n4196;
  LPM_q_ivl_33979 <= tmp_ivl_33981 & tmp_ivl_33976;
  tmp_ivl_33983 <= tmp_ivl_33987(1);
  tmp_ivl_33985 <= tmp_ivl_33987(0);
  tmp_ivl_33987 <= LPM_d0_ivl_33991(0 + 1 downto 0);
  tmp_ivl_33992 <= new_AGEMA_signal_3458 & n4212;
  LPM_q_ivl_33995 <= tmp_ivl_33997 & tmp_ivl_33992;
  tmp_ivl_33999 <= new_AGEMA_signal_3454 & n4213;
  LPM_q_ivl_34002 <= tmp_ivl_34004 & tmp_ivl_33999;
  new_AGEMA_signal_3878 <= tmp_ivl_34006(1);
  n4197 <= tmp_ivl_34006(0);
  tmp_ivl_34006 <= LPM_d0_ivl_34010(0 + 1 downto 0);
  tmp_ivl_34011 <= new_AGEMA_signal_3472 & n4198;
  LPM_q_ivl_34014 <= tmp_ivl_34016 & tmp_ivl_34011;
  tmp_ivl_34018 <= new_AGEMA_signal_3878 & n4197;
  LPM_q_ivl_34021 <= tmp_ivl_34023 & tmp_ivl_34018;
  tmp_ivl_34025 <= tmp_ivl_34029(1);
  tmp_ivl_34027 <= tmp_ivl_34029(0);
  tmp_ivl_34029 <= LPM_d0_ivl_34033(0 + 1 downto 0);
  tmp_ivl_34034 <= new_AGEMA_signal_3469 & n4199;
  LPM_q_ivl_34037 <= tmp_ivl_34039 & tmp_ivl_34034;
  tmp_ivl_34041 <= new_AGEMA_signal_3454 & n4213;
  LPM_q_ivl_34044 <= tmp_ivl_34046 & tmp_ivl_34041;
  new_AGEMA_signal_3879 <= tmp_ivl_34048(1);
  n4200 <= tmp_ivl_34048(0);
  tmp_ivl_34048 <= LPM_d0_ivl_34052(0 + 1 downto 0);
  tmp_ivl_34053 <= new_AGEMA_signal_3879 & n4200;
  LPM_q_ivl_34056 <= tmp_ivl_34058 & tmp_ivl_34053;
  tmp_ivl_34060 <= new_AGEMA_signal_3507 & n4202;
  LPM_q_ivl_34063 <= tmp_ivl_34065 & tmp_ivl_34060;
  tmp_ivl_34067 <= tmp_ivl_34071(1);
  tmp_ivl_34069 <= tmp_ivl_34071(0);
  tmp_ivl_34071 <= LPM_d0_ivl_34075(0 + 1 downto 0);
  tmp_ivl_34076 <= new_AGEMA_signal_4565 & n4219;
  LPM_q_ivl_34079 <= tmp_ivl_34081 & tmp_ivl_34076;
  tmp_ivl_34083 <= new_AGEMA_signal_3467 & n4201;
  LPM_q_ivl_34086 <= tmp_ivl_34088 & tmp_ivl_34083;
  new_AGEMA_signal_4607 <= tmp_ivl_34090(1);
  n4203 <= tmp_ivl_34090(0);
  tmp_ivl_34090 <= LPM_d0_ivl_34094(0 + 1 downto 0);
  tmp_ivl_34095 <= new_AGEMA_signal_4607 & n4203;
  LPM_q_ivl_34098 <= tmp_ivl_34100 & tmp_ivl_34095;
  tmp_ivl_34102 <= new_AGEMA_signal_3507 & n4202;
  LPM_q_ivl_34105 <= tmp_ivl_34107 & tmp_ivl_34102;
  tmp_ivl_34109 <= tmp_ivl_34113(1);
  tmp_ivl_34111 <= tmp_ivl_34113(0);
  tmp_ivl_34113 <= LPM_d0_ivl_34117(0 + 1 downto 0);
  tmp_ivl_34118 <= new_AGEMA_signal_3460 & n4204;
  LPM_q_ivl_34121 <= tmp_ivl_34123 & tmp_ivl_34118;
  tmp_ivl_34125 <= new_AGEMA_signal_4143 & n4228;
  LPM_q_ivl_34128 <= tmp_ivl_34130 & tmp_ivl_34125;
  new_AGEMA_signal_4436 <= tmp_ivl_34132(1);
  n4207 <= tmp_ivl_34132(0);
  tmp_ivl_34132 <= LPM_d0_ivl_34136(0 + 1 downto 0);
  tmp_ivl_34139 <= tmp_ivl_34137 & n4206;
  LPM_q_ivl_34142 <= tmp_ivl_34144 & tmp_ivl_34139;
  tmp_ivl_34146 <= new_AGEMA_signal_3514 & n4205;
  LPM_q_ivl_34149 <= tmp_ivl_34151 & tmp_ivl_34146;
  new_AGEMA_signal_3880 <= tmp_ivl_34153(1);
  n4237 <= tmp_ivl_34153(0);
  tmp_ivl_34153 <= LPM_d0_ivl_34157(0 + 1 downto 0);
  tmp_ivl_34158 <= new_AGEMA_signal_4436 & n4207;
  LPM_q_ivl_34161 <= tmp_ivl_34163 & tmp_ivl_34158;
  tmp_ivl_34165 <= new_AGEMA_signal_3880 & n4237;
  LPM_q_ivl_34168 <= tmp_ivl_34170 & tmp_ivl_34165;
  tmp_ivl_34172 <= tmp_ivl_34176(1);
  tmp_ivl_34174 <= tmp_ivl_34176(0);
  tmp_ivl_34176 <= LPM_d0_ivl_34180(0 + 1 downto 0);
  tmp_ivl_34181 <= new_AGEMA_signal_2843 & n4208;
  LPM_q_ivl_34184 <= tmp_ivl_34186 & tmp_ivl_34181;
  tmp_ivl_34189 <= z2(4);
  tmp_ivl_34190 <= new_AGEMA_signal_3208 & tmp_ivl_34189;
  LPM_q_ivl_34193 <= tmp_ivl_34195 & tmp_ivl_34190;
  new_AGEMA_signal_3516 <= tmp_ivl_34197(1);
  n4209 <= tmp_ivl_34197(0);
  tmp_ivl_34197 <= LPM_d0_ivl_34201(0 + 1 downto 0);
  tmp_ivl_34202 <= new_AGEMA_signal_3829 & n4210;
  LPM_q_ivl_34205 <= tmp_ivl_34207 & tmp_ivl_34202;
  tmp_ivl_34209 <= new_AGEMA_signal_3516 & n4209;
  LPM_q_ivl_34212 <= tmp_ivl_34214 & tmp_ivl_34209;
  new_AGEMA_signal_4195 <= tmp_ivl_34216(1);
  n4211 <= tmp_ivl_34216(0);
  tmp_ivl_34216 <= LPM_d0_ivl_34220(0 + 1 downto 0);
  tmp_ivl_34221 <= new_AGEMA_signal_3458 & n4212;
  LPM_q_ivl_34224 <= tmp_ivl_34226 & tmp_ivl_34221;
  tmp_ivl_34228 <= new_AGEMA_signal_4195 & n4211;
  LPM_q_ivl_34231 <= tmp_ivl_34233 & tmp_ivl_34228;
  tmp_ivl_34235 <= tmp_ivl_34239(1);
  tmp_ivl_34237 <= tmp_ivl_34239(0);
  tmp_ivl_34239 <= LPM_d0_ivl_34243(0 + 1 downto 0);
  tmp_ivl_34244 <= new_AGEMA_signal_4564 & n4262;
  LPM_q_ivl_34247 <= tmp_ivl_34249 & tmp_ivl_34244;
  tmp_ivl_34251 <= new_AGEMA_signal_3454 & n4213;
  LPM_q_ivl_34254 <= tmp_ivl_34256 & tmp_ivl_34251;
  new_AGEMA_signal_4608 <= tmp_ivl_34258(1);
  n4214 <= tmp_ivl_34258(0);
  tmp_ivl_34258 <= LPM_d0_ivl_34262(0 + 1 downto 0);
  tmp_ivl_34263 <= new_AGEMA_signal_4608 & n4214;
  LPM_q_ivl_34266 <= tmp_ivl_34268 & tmp_ivl_34263;
  tmp_ivl_34270 <= new_AGEMA_signal_3510 & n4250;
  LPM_q_ivl_34273 <= tmp_ivl_34275 & tmp_ivl_34270;
  tmp_ivl_34277 <= tmp_ivl_34281(1);
  tmp_ivl_34279 <= tmp_ivl_34281(0);
  tmp_ivl_34281 <= LPM_d0_ivl_34285(0 + 1 downto 0);
  tmp_ivl_34286 <= new_AGEMA_signal_3508 & n4215;
  LPM_q_ivl_34289 <= tmp_ivl_34291 & tmp_ivl_34286;
  tmp_ivl_34293 <= new_AGEMA_signal_3505 & n4220;
  LPM_q_ivl_34296 <= tmp_ivl_34298 & tmp_ivl_34293;
  new_AGEMA_signal_3881 <= tmp_ivl_34300(1);
  n4216 <= tmp_ivl_34300(0);
  tmp_ivl_34300 <= LPM_d0_ivl_34304(0 + 1 downto 0);
  tmp_ivl_34305 <= new_AGEMA_signal_3881 & n4216;
  LPM_q_ivl_34308 <= tmp_ivl_34310 & tmp_ivl_34305;
  tmp_ivl_34312 <= new_AGEMA_signal_4138 & n4217;
  LPM_q_ivl_34315 <= tmp_ivl_34317 & tmp_ivl_34312;
  tmp_ivl_34319 <= tmp_ivl_34323(1);
  tmp_ivl_34321 <= tmp_ivl_34323(0);
  tmp_ivl_34323 <= LPM_d0_ivl_34327(0 + 1 downto 0);
  tmp_ivl_34328 <= new_AGEMA_signal_4138 & n4217;
  LPM_q_ivl_34331 <= tmp_ivl_34333 & tmp_ivl_34328;
  tmp_ivl_34335 <= new_AGEMA_signal_3823 & n4222;
  LPM_q_ivl_34338 <= tmp_ivl_34340 & tmp_ivl_34335;
  new_AGEMA_signal_4439 <= tmp_ivl_34342(1);
  n4218 <= tmp_ivl_34342(0);
  tmp_ivl_34342 <= LPM_d0_ivl_34346(0 + 1 downto 0);
  tmp_ivl_34347 <= new_AGEMA_signal_4565 & n4219;
  LPM_q_ivl_34350 <= tmp_ivl_34352 & tmp_ivl_34347;
  tmp_ivl_34354 <= new_AGEMA_signal_4439 & n4218;
  LPM_q_ivl_34357 <= tmp_ivl_34359 & tmp_ivl_34354;
  tmp_ivl_34361 <= tmp_ivl_34365(1);
  tmp_ivl_34363 <= tmp_ivl_34365(0);
  tmp_ivl_34365 <= LPM_d0_ivl_34369(0 + 1 downto 0);
  tmp_ivl_34370 <= new_AGEMA_signal_3505 & n4220;
  LPM_q_ivl_34373 <= tmp_ivl_34375 & tmp_ivl_34370;
  tmp_ivl_34377 <= new_AGEMA_signal_3504 & n4223;
  LPM_q_ivl_34380 <= tmp_ivl_34382 & tmp_ivl_34377;
  new_AGEMA_signal_3882 <= tmp_ivl_34384(1);
  n4221 <= tmp_ivl_34384(0);
  tmp_ivl_34384 <= LPM_d0_ivl_34388(0 + 1 downto 0);
  tmp_ivl_34389 <= new_AGEMA_signal_3823 & n4222;
  LPM_q_ivl_34392 <= tmp_ivl_34394 & tmp_ivl_34389;
  tmp_ivl_34396 <= new_AGEMA_signal_3882 & n4221;
  LPM_q_ivl_34399 <= tmp_ivl_34401 & tmp_ivl_34396;
  tmp_ivl_34403 <= tmp_ivl_34407(1);
  tmp_ivl_34405 <= tmp_ivl_34407(0);
  tmp_ivl_34407 <= LPM_d0_ivl_34411(0 + 1 downto 0);
  tmp_ivl_34412 <= new_AGEMA_signal_3817 & n4224;
  LPM_q_ivl_34415 <= tmp_ivl_34417 & tmp_ivl_34412;
  tmp_ivl_34419 <= new_AGEMA_signal_3504 & n4223;
  LPM_q_ivl_34422 <= tmp_ivl_34424 & tmp_ivl_34419;
  new_AGEMA_signal_4197 <= tmp_ivl_34426(1);
  n4225 <= tmp_ivl_34426(0);
  tmp_ivl_34426 <= LPM_d0_ivl_34430(0 + 1 downto 0);
  tmp_ivl_34431 <= new_AGEMA_signal_3503 & n4226;
  LPM_q_ivl_34434 <= tmp_ivl_34436 & tmp_ivl_34431;
  tmp_ivl_34438 <= new_AGEMA_signal_4197 & n4225;
  LPM_q_ivl_34441 <= tmp_ivl_34443 & tmp_ivl_34438;
  tmp_ivl_34445 <= tmp_ivl_34449(1);
  tmp_ivl_34447 <= tmp_ivl_34449(0);
  tmp_ivl_34449 <= LPM_d0_ivl_34453(0 + 1 downto 0);
  tmp_ivl_34455 <= z3(6);
  tmp_ivl_34456 <= new_AGEMA_signal_3579 & tmp_ivl_34455;
  LPM_q_ivl_34459 <= tmp_ivl_34461 & tmp_ivl_34456;
  tmp_ivl_34464 <= state_in_s1(254);
  tmp_ivl_34466 <= state_in_s0(254);
  tmp_ivl_34467 <= tmp_ivl_34464 & tmp_ivl_34466;
  LPM_q_ivl_34470 <= tmp_ivl_34472 & tmp_ivl_34467;
  new_AGEMA_signal_3883 <= tmp_ivl_34474(1);
  n4227 <= tmp_ivl_34474(0);
  tmp_ivl_34474 <= LPM_d0_ivl_34478(0 + 1 downto 0);
  tmp_ivl_34479 <= new_AGEMA_signal_4143 & n4228;
  LPM_q_ivl_34482 <= tmp_ivl_34484 & tmp_ivl_34479;
  tmp_ivl_34486 <= new_AGEMA_signal_3883 & n4227;
  LPM_q_ivl_34489 <= tmp_ivl_34491 & tmp_ivl_34486;
  new_AGEMA_signal_4441 <= tmp_ivl_34493(1);
  n4235 <= tmp_ivl_34493(0);
  tmp_ivl_34493 <= LPM_d0_ivl_34497(0 + 1 downto 0);
  tmp_ivl_34498 <= new_AGEMA_signal_4091 & n4230;
  LPM_q_ivl_34501 <= tmp_ivl_34503 & tmp_ivl_34498;
  tmp_ivl_34505 <= new_AGEMA_signal_4100 & n4229;
  LPM_q_ivl_34508 <= tmp_ivl_34510 & tmp_ivl_34505;
  new_AGEMA_signal_4442 <= tmp_ivl_34512(1);
  n4231 <= tmp_ivl_34512(0);
  tmp_ivl_34512 <= LPM_d0_ivl_34516(0 + 1 downto 0);
  tmp_ivl_34517 <= new_AGEMA_signal_4441 & n4235;
  LPM_q_ivl_34520 <= tmp_ivl_34522 & tmp_ivl_34517;
  tmp_ivl_34524 <= new_AGEMA_signal_4442 & n4231;
  LPM_q_ivl_34527 <= tmp_ivl_34529 & tmp_ivl_34524;
  tmp_ivl_34531 <= tmp_ivl_34535(1);
  tmp_ivl_34533 <= tmp_ivl_34535(0);
  tmp_ivl_34535 <= LPM_d0_ivl_34539(0 + 1 downto 0);
  tmp_ivl_34540 <= new_AGEMA_signal_4123 & n4233;
  LPM_q_ivl_34543 <= tmp_ivl_34545 & tmp_ivl_34540;
  tmp_ivl_34547 <= new_AGEMA_signal_4136 & n4232;
  LPM_q_ivl_34550 <= tmp_ivl_34552 & tmp_ivl_34547;
  new_AGEMA_signal_4443 <= tmp_ivl_34554(1);
  n4234 <= tmp_ivl_34554(0);
  tmp_ivl_34554 <= LPM_d0_ivl_34558(0 + 1 downto 0);
  tmp_ivl_34559 <= new_AGEMA_signal_4441 & n4235;
  LPM_q_ivl_34562 <= tmp_ivl_34564 & tmp_ivl_34559;
  tmp_ivl_34566 <= new_AGEMA_signal_4443 & n4234;
  LPM_q_ivl_34569 <= tmp_ivl_34571 & tmp_ivl_34566;
  tmp_ivl_34573 <= tmp_ivl_34577(1);
  tmp_ivl_34575 <= tmp_ivl_34577(0);
  tmp_ivl_34577 <= LPM_d0_ivl_34581(0 + 1 downto 0);
  tmp_ivl_34582 <= new_AGEMA_signal_4441 & n4235;
  LPM_q_ivl_34585 <= tmp_ivl_34587 & tmp_ivl_34582;
  tmp_ivl_34589 <= new_AGEMA_signal_4092 & n4263;
  LPM_q_ivl_34592 <= tmp_ivl_34594 & tmp_ivl_34589;
  new_AGEMA_signal_4570 <= tmp_ivl_34596(1);
  n4236 <= tmp_ivl_34596(0);
  tmp_ivl_34596 <= LPM_d0_ivl_34600(0 + 1 downto 0);
  tmp_ivl_34601 <= new_AGEMA_signal_4570 & n4236;
  LPM_q_ivl_34604 <= tmp_ivl_34606 & tmp_ivl_34601;
  tmp_ivl_34608 <= new_AGEMA_signal_4130 & n4266;
  LPM_q_ivl_34611 <= tmp_ivl_34613 & tmp_ivl_34608;
  tmp_ivl_34615 <= tmp_ivl_34619(1);
  tmp_ivl_34617 <= tmp_ivl_34619(0);
  tmp_ivl_34619 <= LPM_d0_ivl_34623(0 + 1 downto 0);
  tmp_ivl_34625 <= z3(5);
  tmp_ivl_34626 <= new_AGEMA_signal_3574 & tmp_ivl_34625;
  LPM_q_ivl_34629 <= tmp_ivl_34631 & tmp_ivl_34626;
  tmp_ivl_34634 <= state_in_s1(253);
  tmp_ivl_34636 <= state_in_s0(253);
  tmp_ivl_34637 <= tmp_ivl_34634 & tmp_ivl_34636;
  LPM_q_ivl_34640 <= tmp_ivl_34642 & tmp_ivl_34637;
  new_AGEMA_signal_3884 <= tmp_ivl_34644(1);
  n4238 <= tmp_ivl_34644(0);
  tmp_ivl_34644 <= LPM_d0_ivl_34648(0 + 1 downto 0);
  tmp_ivl_34649 <= new_AGEMA_signal_3884 & n4238;
  LPM_q_ivl_34652 <= tmp_ivl_34654 & tmp_ivl_34649;
  tmp_ivl_34656 <= new_AGEMA_signal_3880 & n4237;
  LPM_q_ivl_34659 <= tmp_ivl_34661 & tmp_ivl_34656;
  new_AGEMA_signal_4198 <= tmp_ivl_34663(1);
  n4247 <= tmp_ivl_34663(0);
  tmp_ivl_34663 <= LPM_d0_ivl_34667(0 + 1 downto 0);
  tmp_ivl_34668 <= new_AGEMA_signal_4097 & n4239;
  LPM_q_ivl_34671 <= tmp_ivl_34673 & tmp_ivl_34668;
  tmp_ivl_34675 <= new_AGEMA_signal_4198 & n4247;
  LPM_q_ivl_34678 <= tmp_ivl_34680 & tmp_ivl_34675;
  new_AGEMA_signal_4444 <= tmp_ivl_34682(1);
  n4240 <= tmp_ivl_34682(0);
  tmp_ivl_34682 <= LPM_d0_ivl_34686(0 + 1 downto 0);
  tmp_ivl_34687 <= new_AGEMA_signal_4089 & n4241;
  LPM_q_ivl_34690 <= tmp_ivl_34692 & tmp_ivl_34687;
  tmp_ivl_34694 <= new_AGEMA_signal_4444 & n4240;
  LPM_q_ivl_34697 <= tmp_ivl_34699 & tmp_ivl_34694;
  tmp_ivl_34701 <= tmp_ivl_34705(1);
  tmp_ivl_34703 <= tmp_ivl_34705(0);
  tmp_ivl_34705 <= LPM_d0_ivl_34709(0 + 1 downto 0);
  tmp_ivl_34710 <= new_AGEMA_signal_4122 & n4243;
  LPM_q_ivl_34713 <= tmp_ivl_34715 & tmp_ivl_34710;
  tmp_ivl_34717 <= new_AGEMA_signal_4134 & n4242;
  LPM_q_ivl_34720 <= tmp_ivl_34722 & tmp_ivl_34717;
  new_AGEMA_signal_4445 <= tmp_ivl_34724(1);
  n4244 <= tmp_ivl_34724(0);
  tmp_ivl_34724 <= LPM_d0_ivl_34728(0 + 1 downto 0);
  tmp_ivl_34729 <= new_AGEMA_signal_4445 & n4244;
  LPM_q_ivl_34732 <= tmp_ivl_34734 & tmp_ivl_34729;
  tmp_ivl_34736 <= new_AGEMA_signal_4198 & n4247;
  LPM_q_ivl_34739 <= tmp_ivl_34741 & tmp_ivl_34736;
  tmp_ivl_34743 <= tmp_ivl_34747(1);
  tmp_ivl_34745 <= tmp_ivl_34747(0);
  tmp_ivl_34747 <= LPM_d0_ivl_34751(0 + 1 downto 0);
  tmp_ivl_34752 <= new_AGEMA_signal_4129 & n4246;
  LPM_q_ivl_34755 <= tmp_ivl_34757 & tmp_ivl_34752;
  tmp_ivl_34759 <= new_AGEMA_signal_4088 & n4245;
  LPM_q_ivl_34762 <= tmp_ivl_34764 & tmp_ivl_34759;
  new_AGEMA_signal_4446 <= tmp_ivl_34766(1);
  n4248 <= tmp_ivl_34766(0);
  tmp_ivl_34766 <= LPM_d0_ivl_34770(0 + 1 downto 0);
  tmp_ivl_34771 <= new_AGEMA_signal_4446 & n4248;
  LPM_q_ivl_34774 <= tmp_ivl_34776 & tmp_ivl_34771;
  tmp_ivl_34778 <= new_AGEMA_signal_4198 & n4247;
  LPM_q_ivl_34781 <= tmp_ivl_34783 & tmp_ivl_34778;
  tmp_ivl_34785 <= tmp_ivl_34789(1);
  tmp_ivl_34787 <= tmp_ivl_34789(0);
  tmp_ivl_34789 <= LPM_d0_ivl_34793(0 + 1 downto 0);
  tmp_ivl_34795 <= z3(4);
  tmp_ivl_34796 <= new_AGEMA_signal_3563 & tmp_ivl_34795;
  LPM_q_ivl_34799 <= tmp_ivl_34801 & tmp_ivl_34796;
  tmp_ivl_34804 <= state_in_s1(252);
  tmp_ivl_34806 <= state_in_s0(252);
  tmp_ivl_34807 <= tmp_ivl_34804 & tmp_ivl_34806;
  LPM_q_ivl_34810 <= tmp_ivl_34812 & tmp_ivl_34807;
  new_AGEMA_signal_3885 <= tmp_ivl_34814(1);
  n4249 <= tmp_ivl_34814(0);
  tmp_ivl_34814 <= LPM_d0_ivl_34818(0 + 1 downto 0);
  tmp_ivl_34819 <= new_AGEMA_signal_3510 & n4250;
  LPM_q_ivl_34822 <= tmp_ivl_34824 & tmp_ivl_34819;
  tmp_ivl_34826 <= new_AGEMA_signal_3885 & n4249;
  LPM_q_ivl_34829 <= tmp_ivl_34831 & tmp_ivl_34826;
  new_AGEMA_signal_4199 <= tmp_ivl_34833(1);
  n4260 <= tmp_ivl_34833(0);
  tmp_ivl_34833 <= LPM_d0_ivl_34837(0 + 1 downto 0);
  tmp_ivl_34838 <= new_AGEMA_signal_4199 & n4260;
  LPM_q_ivl_34841 <= tmp_ivl_34843 & tmp_ivl_34838;
  tmp_ivl_34845 <= new_AGEMA_signal_4121 & n4251;
  LPM_q_ivl_34848 <= tmp_ivl_34850 & tmp_ivl_34845;
  new_AGEMA_signal_4447 <= tmp_ivl_34852(1);
  n4252 <= tmp_ivl_34852(0);
  tmp_ivl_34852 <= LPM_d0_ivl_34856(0 + 1 downto 0);
  tmp_ivl_34857 <= new_AGEMA_signal_4133 & n4253;
  LPM_q_ivl_34860 <= tmp_ivl_34862 & tmp_ivl_34857;
  tmp_ivl_34864 <= new_AGEMA_signal_4447 & n4252;
  LPM_q_ivl_34867 <= tmp_ivl_34869 & tmp_ivl_34864;
  tmp_ivl_34871 <= tmp_ivl_34875(1);
  tmp_ivl_34873 <= tmp_ivl_34875(0);
  tmp_ivl_34875 <= LPM_d0_ivl_34879(0 + 1 downto 0);
  tmp_ivl_34880 <= new_AGEMA_signal_4094 & n4255;
  LPM_q_ivl_34883 <= tmp_ivl_34885 & tmp_ivl_34880;
  tmp_ivl_34887 <= new_AGEMA_signal_4086 & n4254;
  LPM_q_ivl_34890 <= tmp_ivl_34892 & tmp_ivl_34887;
  new_AGEMA_signal_4448 <= tmp_ivl_34894(1);
  n4256 <= tmp_ivl_34894(0);
  tmp_ivl_34894 <= LPM_d0_ivl_34898(0 + 1 downto 0);
  tmp_ivl_34899 <= new_AGEMA_signal_4199 & n4260;
  LPM_q_ivl_34902 <= tmp_ivl_34904 & tmp_ivl_34899;
  tmp_ivl_34906 <= new_AGEMA_signal_4448 & n4256;
  LPM_q_ivl_34909 <= tmp_ivl_34911 & tmp_ivl_34906;
  tmp_ivl_34913 <= tmp_ivl_34917(1);
  tmp_ivl_34915 <= tmp_ivl_34917(0);
  tmp_ivl_34917 <= LPM_d0_ivl_34921(0 + 1 downto 0);
  tmp_ivl_34922 <= new_AGEMA_signal_4085 & n4258;
  LPM_q_ivl_34925 <= tmp_ivl_34927 & tmp_ivl_34922;
  tmp_ivl_34929 <= new_AGEMA_signal_4128 & n4257;
  LPM_q_ivl_34932 <= tmp_ivl_34934 & tmp_ivl_34929;
  new_AGEMA_signal_4449 <= tmp_ivl_34936(1);
  n4259 <= tmp_ivl_34936(0);
  tmp_ivl_34936 <= LPM_d0_ivl_34940(0 + 1 downto 0);
  tmp_ivl_34941 <= new_AGEMA_signal_4199 & n4260;
  LPM_q_ivl_34944 <= tmp_ivl_34946 & tmp_ivl_34941;
  tmp_ivl_34948 <= new_AGEMA_signal_4449 & n4259;
  LPM_q_ivl_34951 <= tmp_ivl_34953 & tmp_ivl_34948;
  tmp_ivl_34955 <= tmp_ivl_34959(1);
  tmp_ivl_34957 <= tmp_ivl_34959(0);
  tmp_ivl_34959 <= LPM_d0_ivl_34963(0 + 1 downto 0);
  tmp_ivl_34965 <= z3(3);
  tmp_ivl_34966 <= new_AGEMA_signal_3552 & tmp_ivl_34965;
  LPM_q_ivl_34969 <= tmp_ivl_34971 & tmp_ivl_34966;
  tmp_ivl_34974 <= state_in_s1(251);
  tmp_ivl_34976 <= state_in_s0(251);
  tmp_ivl_34977 <= tmp_ivl_34974 & tmp_ivl_34976;
  LPM_q_ivl_34980 <= tmp_ivl_34982 & tmp_ivl_34977;
  new_AGEMA_signal_3886 <= tmp_ivl_34984(1);
  n4261 <= tmp_ivl_34984(0);
  tmp_ivl_34984 <= LPM_d0_ivl_34988(0 + 1 downto 0);
  tmp_ivl_34989 <= new_AGEMA_signal_4564 & n4262;
  LPM_q_ivl_34992 <= tmp_ivl_34994 & tmp_ivl_34989;
  tmp_ivl_34996 <= new_AGEMA_signal_3886 & n4261;
  LPM_q_ivl_34999 <= tmp_ivl_35001 & tmp_ivl_34996;
  new_AGEMA_signal_4611 <= tmp_ivl_35003(1);
  n4272 <= tmp_ivl_35003(0);
  tmp_ivl_35003 <= LPM_d0_ivl_35007(0 + 1 downto 0);
  tmp_ivl_35008 <= new_AGEMA_signal_4082 & n4264;
  LPM_q_ivl_35011 <= tmp_ivl_35013 & tmp_ivl_35008;
  tmp_ivl_35015 <= new_AGEMA_signal_4092 & n4263;
  LPM_q_ivl_35018 <= tmp_ivl_35020 & tmp_ivl_35015;
  new_AGEMA_signal_4450 <= tmp_ivl_35022(1);
  n4265 <= tmp_ivl_35022(0);
  tmp_ivl_35022 <= LPM_d0_ivl_35026(0 + 1 downto 0);
  tmp_ivl_35027 <= new_AGEMA_signal_4611 & n4272;
  LPM_q_ivl_35030 <= tmp_ivl_35032 & tmp_ivl_35027;
  tmp_ivl_35034 <= new_AGEMA_signal_4450 & n4265;
  LPM_q_ivl_35037 <= tmp_ivl_35039 & tmp_ivl_35034;
  tmp_ivl_35041 <= tmp_ivl_35045(1);
  tmp_ivl_35043 <= tmp_ivl_35045(0);
  tmp_ivl_35045 <= LPM_d0_ivl_35049(0 + 1 downto 0);
  tmp_ivl_35050 <= new_AGEMA_signal_4120 & n4267;
  LPM_q_ivl_35053 <= tmp_ivl_35055 & tmp_ivl_35050;
  tmp_ivl_35057 <= new_AGEMA_signal_4130 & n4266;
  LPM_q_ivl_35060 <= tmp_ivl_35062 & tmp_ivl_35057;
  new_AGEMA_signal_4451 <= tmp_ivl_35064(1);
  n4268 <= tmp_ivl_35064(0);
  tmp_ivl_35064 <= LPM_d0_ivl_35068(0 + 1 downto 0);
  tmp_ivl_35069 <= new_AGEMA_signal_4611 & n4272;
  LPM_q_ivl_35072 <= tmp_ivl_35074 & tmp_ivl_35069;
  tmp_ivl_35076 <= new_AGEMA_signal_4451 & n4268;
  LPM_q_ivl_35079 <= tmp_ivl_35081 & tmp_ivl_35076;
  tmp_ivl_35083 <= tmp_ivl_35087(1);
  tmp_ivl_35085 <= tmp_ivl_35087(0);
  tmp_ivl_35087 <= LPM_d0_ivl_35091(0 + 1 downto 0);
  tmp_ivl_35092 <= new_AGEMA_signal_4127 & n4270;
  LPM_q_ivl_35095 <= tmp_ivl_35097 & tmp_ivl_35092;
  tmp_ivl_35099 <= new_AGEMA_signal_4083 & n4269;
  LPM_q_ivl_35102 <= tmp_ivl_35104 & tmp_ivl_35099;
  new_AGEMA_signal_4452 <= tmp_ivl_35106(1);
  n4271 <= tmp_ivl_35106(0);
  tmp_ivl_35106 <= LPM_d0_ivl_35110(0 + 1 downto 0);
  tmp_ivl_35111 <= new_AGEMA_signal_4611 & n4272;
  LPM_q_ivl_35114 <= tmp_ivl_35116 & tmp_ivl_35111;
  tmp_ivl_35118 <= new_AGEMA_signal_4452 & n4271;
  LPM_q_ivl_35121 <= tmp_ivl_35123 & tmp_ivl_35118;
  tmp_ivl_35125 <= tmp_ivl_35129(1);
  tmp_ivl_35127 <= tmp_ivl_35129(0);
  tmp_ivl_35129 <= LPM_d0_ivl_35133(0 + 1 downto 0);
  tmp_ivl_35135 <= y2(0);
  tmp_ivl_35136 <= new_AGEMA_signal_2989 & tmp_ivl_35135;
  LPM_q_ivl_35139 <= tmp_ivl_35141 & tmp_ivl_35136;
  tmp_ivl_35143 <= new_AGEMA_signal_2890 & SboxInst_n384;
  LPM_q_ivl_35146 <= tmp_ivl_35148 & tmp_ivl_35143;
  tmp_ivl_35151 <= fresh(0);
  LPM_q_ivl_35153 <= tmp_ivl_35155 & tmp_ivl_35151;
  new_AGEMA_signal_3517 <= tmp_ivl_35159(1);
  tmp_ivl_35157 <= tmp_ivl_35159(0);
  tmp_ivl_35159 <= LPM_d0_ivl_35163(0 + 1 downto 0);
  tmp_ivl_35164 <= new_AGEMA_signal_2704 & n3290;
  LPM_q_ivl_35167 <= tmp_ivl_35169 & tmp_ivl_35164;
  tmp_ivl_35171 <= new_AGEMA_signal_2979 & SboxInst_n383;
  LPM_q_ivl_35174 <= tmp_ivl_35176 & tmp_ivl_35171;
  tmp_ivl_35179 <= fresh(1);
  LPM_q_ivl_35181 <= tmp_ivl_35183 & tmp_ivl_35179;
  new_AGEMA_signal_2991 <= tmp_ivl_35187(1);
  tmp_ivl_35185 <= tmp_ivl_35187(0);
  tmp_ivl_35187 <= LPM_d0_ivl_35191(0 + 1 downto 0);
  tmp_ivl_35192 <= new_AGEMA_signal_2709 & n3289;
  LPM_q_ivl_35195 <= tmp_ivl_35197 & tmp_ivl_35192;
  tmp_ivl_35199 <= new_AGEMA_signal_2977 & SboxInst_n382;
  LPM_q_ivl_35202 <= tmp_ivl_35204 & tmp_ivl_35199;
  tmp_ivl_35207 <= fresh(2);
  LPM_q_ivl_35209 <= tmp_ivl_35211 & tmp_ivl_35207;
  new_AGEMA_signal_2992 <= tmp_ivl_35215(1);
  tmp_ivl_35213 <= tmp_ivl_35215(0);
  tmp_ivl_35215 <= LPM_d0_ivl_35219(0 + 1 downto 0);
  tmp_ivl_35220 <= new_AGEMA_signal_2717 & n3288;
  LPM_q_ivl_35223 <= tmp_ivl_35225 & tmp_ivl_35220;
  tmp_ivl_35227 <= new_AGEMA_signal_2975 & SboxInst_n381;
  LPM_q_ivl_35230 <= tmp_ivl_35232 & tmp_ivl_35227;
  tmp_ivl_35235 <= fresh(3);
  LPM_q_ivl_35237 <= tmp_ivl_35239 & tmp_ivl_35235;
  new_AGEMA_signal_2993 <= tmp_ivl_35243(1);
  tmp_ivl_35241 <= tmp_ivl_35243(0);
  tmp_ivl_35243 <= LPM_d0_ivl_35247(0 + 1 downto 0);
  tmp_ivl_35248 <= new_AGEMA_signal_2727 & n3286;
  LPM_q_ivl_35251 <= tmp_ivl_35253 & tmp_ivl_35248;
  tmp_ivl_35255 <= new_AGEMA_signal_2974 & SboxInst_n380;
  LPM_q_ivl_35258 <= tmp_ivl_35260 & tmp_ivl_35255;
  tmp_ivl_35263 <= fresh(4);
  LPM_q_ivl_35265 <= tmp_ivl_35267 & tmp_ivl_35263;
  new_AGEMA_signal_2994 <= tmp_ivl_35271(1);
  tmp_ivl_35269 <= tmp_ivl_35271(0);
  tmp_ivl_35271 <= LPM_d0_ivl_35275(0 + 1 downto 0);
  tmp_ivl_35276 <= new_AGEMA_signal_2733 & n3285;
  LPM_q_ivl_35279 <= tmp_ivl_35281 & tmp_ivl_35276;
  tmp_ivl_35283 <= new_AGEMA_signal_2971 & SboxInst_n379;
  LPM_q_ivl_35286 <= tmp_ivl_35288 & tmp_ivl_35283;
  tmp_ivl_35291 <= fresh(5);
  LPM_q_ivl_35293 <= tmp_ivl_35295 & tmp_ivl_35291;
  new_AGEMA_signal_2995 <= tmp_ivl_35299(1);
  tmp_ivl_35297 <= tmp_ivl_35299(0);
  tmp_ivl_35299 <= LPM_d0_ivl_35303(0 + 1 downto 0);
  tmp_ivl_35304 <= new_AGEMA_signal_2742 & n3284;
  LPM_q_ivl_35307 <= tmp_ivl_35309 & tmp_ivl_35304;
  tmp_ivl_35311 <= new_AGEMA_signal_2970 & SboxInst_n378;
  LPM_q_ivl_35314 <= tmp_ivl_35316 & tmp_ivl_35311;
  tmp_ivl_35319 <= fresh(6);
  LPM_q_ivl_35321 <= tmp_ivl_35323 & tmp_ivl_35319;
  new_AGEMA_signal_2996 <= tmp_ivl_35327(1);
  tmp_ivl_35325 <= tmp_ivl_35327(0);
  tmp_ivl_35327 <= LPM_d0_ivl_35331(0 + 1 downto 0);
  tmp_ivl_35332 <= new_AGEMA_signal_2750 & n3283;
  LPM_q_ivl_35335 <= tmp_ivl_35337 & tmp_ivl_35332;
  tmp_ivl_35339 <= new_AGEMA_signal_2968 & SboxInst_n377;
  LPM_q_ivl_35342 <= tmp_ivl_35344 & tmp_ivl_35339;
  tmp_ivl_35347 <= fresh(7);
  LPM_q_ivl_35349 <= tmp_ivl_35351 & tmp_ivl_35347;
  new_AGEMA_signal_2997 <= tmp_ivl_35355(1);
  tmp_ivl_35353 <= tmp_ivl_35355(0);
  tmp_ivl_35355 <= LPM_d0_ivl_35359(0 + 1 downto 0);
  tmp_ivl_35360 <= new_AGEMA_signal_2755 & n3282;
  LPM_q_ivl_35363 <= tmp_ivl_35365 & tmp_ivl_35360;
  tmp_ivl_35367 <= new_AGEMA_signal_2964 & SboxInst_n376;
  LPM_q_ivl_35370 <= tmp_ivl_35372 & tmp_ivl_35367;
  tmp_ivl_35375 <= fresh(8);
  LPM_q_ivl_35377 <= tmp_ivl_35379 & tmp_ivl_35375;
  new_AGEMA_signal_2998 <= tmp_ivl_35383(1);
  tmp_ivl_35381 <= tmp_ivl_35383(0);
  tmp_ivl_35383 <= LPM_d0_ivl_35387(0 + 1 downto 0);
  tmp_ivl_35388 <= new_AGEMA_signal_2760 & n3281;
  LPM_q_ivl_35391 <= tmp_ivl_35393 & tmp_ivl_35388;
  tmp_ivl_35395 <= new_AGEMA_signal_2978 & SboxInst_n375;
  LPM_q_ivl_35398 <= tmp_ivl_35400 & tmp_ivl_35395;
  tmp_ivl_35403 <= fresh(9);
  LPM_q_ivl_35405 <= tmp_ivl_35407 & tmp_ivl_35403;
  new_AGEMA_signal_2999 <= tmp_ivl_35411(1);
  tmp_ivl_35409 <= tmp_ivl_35411(0);
  tmp_ivl_35411 <= LPM_d0_ivl_35415(0 + 1 downto 0);
  tmp_ivl_35416 <= new_AGEMA_signal_2695 & n3280;
  LPM_q_ivl_35419 <= tmp_ivl_35421 & tmp_ivl_35416;
  tmp_ivl_35423 <= new_AGEMA_signal_2976 & SboxInst_n374;
  LPM_q_ivl_35426 <= tmp_ivl_35428 & tmp_ivl_35423;
  tmp_ivl_35431 <= fresh(10);
  LPM_q_ivl_35433 <= tmp_ivl_35435 & tmp_ivl_35431;
  new_AGEMA_signal_3000 <= tmp_ivl_35439(1);
  tmp_ivl_35437 <= tmp_ivl_35439(0);
  tmp_ivl_35439 <= LPM_d0_ivl_35443(0 + 1 downto 0);
  tmp_ivl_35445 <= y2(1);
  tmp_ivl_35446 <= new_AGEMA_signal_3513 & tmp_ivl_35445;
  LPM_q_ivl_35449 <= tmp_ivl_35451 & tmp_ivl_35446;
  tmp_ivl_35453 <= new_AGEMA_signal_2896 & SboxInst_n373;
  LPM_q_ivl_35456 <= tmp_ivl_35458 & tmp_ivl_35453;
  tmp_ivl_35461 <= fresh(11);
  LPM_q_ivl_35463 <= tmp_ivl_35465 & tmp_ivl_35461;
  new_AGEMA_signal_3887 <= tmp_ivl_35469(1);
  tmp_ivl_35467 <= tmp_ivl_35469(0);
  tmp_ivl_35469 <= LPM_d0_ivl_35473(0 + 1 downto 0);
  tmp_ivl_35474 <= new_AGEMA_signal_2701 & n3279;
  LPM_q_ivl_35477 <= tmp_ivl_35479 & tmp_ivl_35474;
  tmp_ivl_35481 <= new_AGEMA_signal_2973 & SboxInst_n372;
  LPM_q_ivl_35484 <= tmp_ivl_35486 & tmp_ivl_35481;
  tmp_ivl_35489 <= fresh(12);
  LPM_q_ivl_35491 <= tmp_ivl_35493 & tmp_ivl_35489;
  new_AGEMA_signal_3001 <= tmp_ivl_35497(1);
  tmp_ivl_35495 <= tmp_ivl_35497(0);
  tmp_ivl_35497 <= LPM_d0_ivl_35501(0 + 1 downto 0);
  tmp_ivl_35502 <= new_AGEMA_signal_2712 & n3278;
  LPM_q_ivl_35505 <= tmp_ivl_35507 & tmp_ivl_35502;
  tmp_ivl_35509 <= new_AGEMA_signal_2972 & SboxInst_n371;
  LPM_q_ivl_35512 <= tmp_ivl_35514 & tmp_ivl_35509;
  tmp_ivl_35517 <= fresh(13);
  LPM_q_ivl_35519 <= tmp_ivl_35521 & tmp_ivl_35517;
  new_AGEMA_signal_3002 <= tmp_ivl_35525(1);
  tmp_ivl_35523 <= tmp_ivl_35525(0);
  tmp_ivl_35525 <= LPM_d0_ivl_35529(0 + 1 downto 0);
  tmp_ivl_35530 <= new_AGEMA_signal_2719 & n3277;
  LPM_q_ivl_35533 <= tmp_ivl_35535 & tmp_ivl_35530;
  tmp_ivl_35537 <= new_AGEMA_signal_2969 & SboxInst_n370;
  LPM_q_ivl_35540 <= tmp_ivl_35542 & tmp_ivl_35537;
  tmp_ivl_35545 <= fresh(14);
  LPM_q_ivl_35547 <= tmp_ivl_35549 & tmp_ivl_35545;
  new_AGEMA_signal_3003 <= tmp_ivl_35553(1);
  tmp_ivl_35551 <= tmp_ivl_35553(0);
  tmp_ivl_35553 <= LPM_d0_ivl_35557(0 + 1 downto 0);
  tmp_ivl_35558 <= new_AGEMA_signal_2724 & n3276;
  LPM_q_ivl_35561 <= tmp_ivl_35563 & tmp_ivl_35558;
  tmp_ivl_35565 <= new_AGEMA_signal_2967 & SboxInst_n369;
  LPM_q_ivl_35568 <= tmp_ivl_35570 & tmp_ivl_35565;
  tmp_ivl_35573 <= fresh(15);
  LPM_q_ivl_35575 <= tmp_ivl_35577 & tmp_ivl_35573;
  new_AGEMA_signal_3004 <= tmp_ivl_35581(1);
  tmp_ivl_35579 <= tmp_ivl_35581(0);
  tmp_ivl_35581 <= LPM_d0_ivl_35585(0 + 1 downto 0);
  tmp_ivl_35586 <= new_AGEMA_signal_2736 & n3275;
  LPM_q_ivl_35589 <= tmp_ivl_35591 & tmp_ivl_35586;
  tmp_ivl_35593 <= new_AGEMA_signal_2965 & SboxInst_n368;
  LPM_q_ivl_35596 <= tmp_ivl_35598 & tmp_ivl_35593;
  tmp_ivl_35601 <= fresh(16);
  LPM_q_ivl_35603 <= tmp_ivl_35605 & tmp_ivl_35601;
  new_AGEMA_signal_3005 <= tmp_ivl_35609(1);
  tmp_ivl_35607 <= tmp_ivl_35609(0);
  tmp_ivl_35609 <= LPM_d0_ivl_35613(0 + 1 downto 0);
  tmp_ivl_35614 <= new_AGEMA_signal_2744 & n3274;
  LPM_q_ivl_35617 <= tmp_ivl_35619 & tmp_ivl_35614;
  tmp_ivl_35621 <= new_AGEMA_signal_2980 & SboxInst_n367;
  LPM_q_ivl_35624 <= tmp_ivl_35626 & tmp_ivl_35621;
  tmp_ivl_35629 <= fresh(17);
  LPM_q_ivl_35631 <= tmp_ivl_35633 & tmp_ivl_35629;
  new_AGEMA_signal_3006 <= tmp_ivl_35637(1);
  tmp_ivl_35635 <= tmp_ivl_35637(0);
  tmp_ivl_35637 <= LPM_d0_ivl_35641(0 + 1 downto 0);
  tmp_ivl_35642 <= new_AGEMA_signal_2698 & n3273;
  LPM_q_ivl_35645 <= tmp_ivl_35647 & tmp_ivl_35642;
  tmp_ivl_35649 <= new_AGEMA_signal_2987 & SboxInst_n366;
  LPM_q_ivl_35652 <= tmp_ivl_35654 & tmp_ivl_35649;
  tmp_ivl_35657 <= fresh(18);
  LPM_q_ivl_35659 <= tmp_ivl_35661 & tmp_ivl_35657;
  new_AGEMA_signal_3007 <= tmp_ivl_35665(1);
  tmp_ivl_35663 <= tmp_ivl_35665(0);
  tmp_ivl_35665 <= LPM_d0_ivl_35669(0 + 1 downto 0);
  tmp_ivl_35670 <= new_AGEMA_signal_2707 & n3272;
  LPM_q_ivl_35673 <= tmp_ivl_35675 & tmp_ivl_35670;
  tmp_ivl_35677 <= new_AGEMA_signal_2985 & SboxInst_n365;
  LPM_q_ivl_35680 <= tmp_ivl_35682 & tmp_ivl_35677;
  tmp_ivl_35685 <= fresh(19);
  LPM_q_ivl_35687 <= tmp_ivl_35689 & tmp_ivl_35685;
  new_AGEMA_signal_3008 <= tmp_ivl_35693(1);
  tmp_ivl_35691 <= tmp_ivl_35693(0);
  tmp_ivl_35693 <= LPM_d0_ivl_35697(0 + 1 downto 0);
  tmp_ivl_35698 <= new_AGEMA_signal_2714 & n3271;
  LPM_q_ivl_35701 <= tmp_ivl_35703 & tmp_ivl_35698;
  tmp_ivl_35705 <= new_AGEMA_signal_2984 & SboxInst_n364;
  LPM_q_ivl_35708 <= tmp_ivl_35710 & tmp_ivl_35705;
  tmp_ivl_35713 <= fresh(20);
  LPM_q_ivl_35715 <= tmp_ivl_35717 & tmp_ivl_35713;
  new_AGEMA_signal_3009 <= tmp_ivl_35721(1);
  tmp_ivl_35719 <= tmp_ivl_35721(0);
  tmp_ivl_35721 <= LPM_d0_ivl_35725(0 + 1 downto 0);
  tmp_ivl_35726 <= new_AGEMA_signal_2721 & n3270;
  LPM_q_ivl_35729 <= tmp_ivl_35731 & tmp_ivl_35726;
  tmp_ivl_35733 <= new_AGEMA_signal_2983 & SboxInst_n363;
  LPM_q_ivl_35736 <= tmp_ivl_35738 & tmp_ivl_35733;
  tmp_ivl_35741 <= fresh(21);
  LPM_q_ivl_35743 <= tmp_ivl_35745 & tmp_ivl_35741;
  new_AGEMA_signal_3010 <= tmp_ivl_35749(1);
  tmp_ivl_35747 <= tmp_ivl_35749(0);
  tmp_ivl_35749 <= LPM_d0_ivl_35753(0 + 1 downto 0);
  tmp_ivl_35754 <= new_AGEMA_signal_3824 & n3287;
  LPM_q_ivl_35757 <= tmp_ivl_35759 & tmp_ivl_35754;
  tmp_ivl_35761 <= new_AGEMA_signal_2895 & SboxInst_n362;
  LPM_q_ivl_35764 <= tmp_ivl_35766 & tmp_ivl_35761;
  tmp_ivl_35769 <= fresh(22);
  LPM_q_ivl_35771 <= tmp_ivl_35773 & tmp_ivl_35769;
  new_AGEMA_signal_4200 <= tmp_ivl_35777(1);
  tmp_ivl_35775 <= tmp_ivl_35777(0);
  tmp_ivl_35777 <= LPM_d0_ivl_35781(0 + 1 downto 0);
  tmp_ivl_35782 <= new_AGEMA_signal_2730 & n3269;
  LPM_q_ivl_35785 <= tmp_ivl_35787 & tmp_ivl_35782;
  tmp_ivl_35789 <= new_AGEMA_signal_2982 & SboxInst_n361;
  LPM_q_ivl_35792 <= tmp_ivl_35794 & tmp_ivl_35789;
  tmp_ivl_35797 <= fresh(23);
  LPM_q_ivl_35799 <= tmp_ivl_35801 & tmp_ivl_35797;
  new_AGEMA_signal_3011 <= tmp_ivl_35805(1);
  tmp_ivl_35803 <= tmp_ivl_35805(0);
  tmp_ivl_35805 <= LPM_d0_ivl_35809(0 + 1 downto 0);
  tmp_ivl_35810 <= new_AGEMA_signal_2739 & n3268;
  LPM_q_ivl_35813 <= tmp_ivl_35815 & tmp_ivl_35810;
  tmp_ivl_35817 <= new_AGEMA_signal_2981 & SboxInst_n360;
  LPM_q_ivl_35820 <= tmp_ivl_35822 & tmp_ivl_35817;
  tmp_ivl_35825 <= fresh(24);
  LPM_q_ivl_35827 <= tmp_ivl_35829 & tmp_ivl_35825;
  new_AGEMA_signal_3012 <= tmp_ivl_35833(1);
  tmp_ivl_35831 <= tmp_ivl_35833(0);
  tmp_ivl_35833 <= LPM_d0_ivl_35837(0 + 1 downto 0);
  tmp_ivl_35838 <= new_AGEMA_signal_2747 & n3267;
  LPM_q_ivl_35841 <= tmp_ivl_35843 & tmp_ivl_35838;
  tmp_ivl_35845 <= new_AGEMA_signal_2872 & SboxInst_n359;
  LPM_q_ivl_35848 <= tmp_ivl_35850 & tmp_ivl_35845;
  tmp_ivl_35853 <= fresh(25);
  LPM_q_ivl_35855 <= tmp_ivl_35857 & tmp_ivl_35853;
  new_AGEMA_signal_3013 <= tmp_ivl_35861(1);
  tmp_ivl_35859 <= tmp_ivl_35861(0);
  tmp_ivl_35861 <= LPM_d0_ivl_35865(0 + 1 downto 0);
  tmp_ivl_35866 <= new_AGEMA_signal_2753 & n3266;
  LPM_q_ivl_35869 <= tmp_ivl_35871 & tmp_ivl_35866;
  tmp_ivl_35873 <= new_AGEMA_signal_2871 & SboxInst_n358;
  LPM_q_ivl_35876 <= tmp_ivl_35878 & tmp_ivl_35873;
  tmp_ivl_35881 <= fresh(26);
  LPM_q_ivl_35883 <= tmp_ivl_35885 & tmp_ivl_35881;
  new_AGEMA_signal_3014 <= tmp_ivl_35889(1);
  tmp_ivl_35887 <= tmp_ivl_35889(0);
  tmp_ivl_35889 <= LPM_d0_ivl_35893(0 + 1 downto 0);
  tmp_ivl_35894 <= new_AGEMA_signal_2758 & n3265;
  LPM_q_ivl_35897 <= tmp_ivl_35899 & tmp_ivl_35894;
  tmp_ivl_35901 <= new_AGEMA_signal_2870 & SboxInst_n357;
  LPM_q_ivl_35904 <= tmp_ivl_35906 & tmp_ivl_35901;
  tmp_ivl_35909 <= fresh(27);
  LPM_q_ivl_35911 <= tmp_ivl_35913 & tmp_ivl_35909;
  new_AGEMA_signal_3015 <= tmp_ivl_35917(1);
  tmp_ivl_35915 <= tmp_ivl_35917(0);
  tmp_ivl_35917 <= LPM_d0_ivl_35921(0 + 1 downto 0);
  tmp_ivl_35922 <= new_AGEMA_signal_2763 & n3264;
  LPM_q_ivl_35925 <= tmp_ivl_35927 & tmp_ivl_35922;
  tmp_ivl_35929 <= new_AGEMA_signal_2869 & SboxInst_n356;
  LPM_q_ivl_35932 <= tmp_ivl_35934 & tmp_ivl_35929;
  tmp_ivl_35937 <= fresh(28);
  LPM_q_ivl_35939 <= tmp_ivl_35941 & tmp_ivl_35937;
  new_AGEMA_signal_3016 <= tmp_ivl_35945(1);
  tmp_ivl_35943 <= tmp_ivl_35945(0);
  tmp_ivl_35945 <= LPM_d0_ivl_35949(0 + 1 downto 0);
  tmp_ivl_35950 <= new_AGEMA_signal_2766 & n3263;
  LPM_q_ivl_35953 <= tmp_ivl_35955 & tmp_ivl_35950;
  tmp_ivl_35957 <= new_AGEMA_signal_2867 & SboxInst_n355;
  LPM_q_ivl_35960 <= tmp_ivl_35962 & tmp_ivl_35957;
  tmp_ivl_35965 <= fresh(29);
  LPM_q_ivl_35967 <= tmp_ivl_35969 & tmp_ivl_35965;
  new_AGEMA_signal_3017 <= tmp_ivl_35973(1);
  tmp_ivl_35971 <= tmp_ivl_35973(0);
  tmp_ivl_35973 <= LPM_d0_ivl_35977(0 + 1 downto 0);
  tmp_ivl_35978 <= new_AGEMA_signal_2769 & n3262;
  LPM_q_ivl_35981 <= tmp_ivl_35983 & tmp_ivl_35978;
  tmp_ivl_35985 <= new_AGEMA_signal_2865 & SboxInst_n354;
  LPM_q_ivl_35988 <= tmp_ivl_35990 & tmp_ivl_35985;
  tmp_ivl_35993 <= fresh(30);
  LPM_q_ivl_35995 <= tmp_ivl_35997 & tmp_ivl_35993;
  new_AGEMA_signal_3018 <= tmp_ivl_36001(1);
  tmp_ivl_35999 <= tmp_ivl_36001(0);
  tmp_ivl_36001 <= LPM_d0_ivl_36005(0 + 1 downto 0);
  tmp_ivl_36006 <= new_AGEMA_signal_2772 & n3261;
  LPM_q_ivl_36009 <= tmp_ivl_36011 & tmp_ivl_36006;
  tmp_ivl_36013 <= new_AGEMA_signal_2863 & SboxInst_n353;
  LPM_q_ivl_36016 <= tmp_ivl_36018 & tmp_ivl_36013;
  tmp_ivl_36021 <= fresh(31);
  LPM_q_ivl_36023 <= tmp_ivl_36025 & tmp_ivl_36021;
  new_AGEMA_signal_3019 <= tmp_ivl_36029(1);
  tmp_ivl_36027 <= tmp_ivl_36029(0);
  tmp_ivl_36029 <= LPM_d0_ivl_36033(0 + 1 downto 0);
  tmp_ivl_36034 <= new_AGEMA_signal_2775 & n3260;
  LPM_q_ivl_36037 <= tmp_ivl_36039 & tmp_ivl_36034;
  tmp_ivl_36041 <= new_AGEMA_signal_2860 & SboxInst_n352;
  LPM_q_ivl_36044 <= tmp_ivl_36046 & tmp_ivl_36041;
  tmp_ivl_36049 <= fresh(32);
  LPM_q_ivl_36051 <= tmp_ivl_36053 & tmp_ivl_36049;
  new_AGEMA_signal_3020 <= tmp_ivl_36057(1);
  tmp_ivl_36055 <= tmp_ivl_36057(0);
  tmp_ivl_36057 <= LPM_d0_ivl_36061(0 + 1 downto 0);
  tmp_ivl_36062 <= new_AGEMA_signal_4432 & n3233;
  LPM_q_ivl_36065 <= tmp_ivl_36067 & tmp_ivl_36062;
  tmp_ivl_36069 <= new_AGEMA_signal_2894 & SboxInst_n351;
  LPM_q_ivl_36072 <= tmp_ivl_36074 & tmp_ivl_36069;
  tmp_ivl_36077 <= fresh(33);
  LPM_q_ivl_36079 <= tmp_ivl_36081 & tmp_ivl_36077;
  new_AGEMA_signal_4577 <= tmp_ivl_36085(1);
  tmp_ivl_36083 <= tmp_ivl_36085(0);
  tmp_ivl_36085 <= LPM_d0_ivl_36089(0 + 1 downto 0);
  tmp_ivl_36090 <= new_AGEMA_signal_2778 & n3259;
  LPM_q_ivl_36093 <= tmp_ivl_36095 & tmp_ivl_36090;
  tmp_ivl_36097 <= new_AGEMA_signal_2861 & SboxInst_n350;
  LPM_q_ivl_36100 <= tmp_ivl_36102 & tmp_ivl_36097;
  tmp_ivl_36105 <= fresh(34);
  LPM_q_ivl_36107 <= tmp_ivl_36109 & tmp_ivl_36105;
  new_AGEMA_signal_3021 <= tmp_ivl_36113(1);
  tmp_ivl_36111 <= tmp_ivl_36113(0);
  tmp_ivl_36113 <= LPM_d0_ivl_36117(0 + 1 downto 0);
  tmp_ivl_36118 <= new_AGEMA_signal_2780 & n3258;
  LPM_q_ivl_36121 <= tmp_ivl_36123 & tmp_ivl_36118;
  tmp_ivl_36125 <= new_AGEMA_signal_2868 & SboxInst_n349;
  LPM_q_ivl_36128 <= tmp_ivl_36130 & tmp_ivl_36125;
  tmp_ivl_36133 <= fresh(35);
  LPM_q_ivl_36135 <= tmp_ivl_36137 & tmp_ivl_36133;
  new_AGEMA_signal_3022 <= tmp_ivl_36141(1);
  tmp_ivl_36139 <= tmp_ivl_36141(0);
  tmp_ivl_36141 <= LPM_d0_ivl_36145(0 + 1 downto 0);
  tmp_ivl_36146 <= new_AGEMA_signal_2783 & n3257;
  LPM_q_ivl_36149 <= tmp_ivl_36151 & tmp_ivl_36146;
  tmp_ivl_36153 <= new_AGEMA_signal_2866 & SboxInst_n348;
  LPM_q_ivl_36156 <= tmp_ivl_36158 & tmp_ivl_36153;
  tmp_ivl_36161 <= fresh(36);
  LPM_q_ivl_36163 <= tmp_ivl_36165 & tmp_ivl_36161;
  new_AGEMA_signal_3023 <= tmp_ivl_36169(1);
  tmp_ivl_36167 <= tmp_ivl_36169(0);
  tmp_ivl_36169 <= LPM_d0_ivl_36173(0 + 1 downto 0);
  tmp_ivl_36174 <= new_AGEMA_signal_2786 & n3256;
  LPM_q_ivl_36177 <= tmp_ivl_36179 & tmp_ivl_36174;
  tmp_ivl_36181 <= new_AGEMA_signal_2864 & SboxInst_n347;
  LPM_q_ivl_36184 <= tmp_ivl_36186 & tmp_ivl_36181;
  tmp_ivl_36189 <= fresh(37);
  LPM_q_ivl_36191 <= tmp_ivl_36193 & tmp_ivl_36189;
  new_AGEMA_signal_3024 <= tmp_ivl_36197(1);
  tmp_ivl_36195 <= tmp_ivl_36197(0);
  tmp_ivl_36197 <= LPM_d0_ivl_36201(0 + 1 downto 0);
  tmp_ivl_36202 <= new_AGEMA_signal_2788 & n3255;
  LPM_q_ivl_36205 <= tmp_ivl_36207 & tmp_ivl_36202;
  tmp_ivl_36209 <= new_AGEMA_signal_2862 & SboxInst_n346;
  LPM_q_ivl_36212 <= tmp_ivl_36214 & tmp_ivl_36209;
  tmp_ivl_36217 <= fresh(38);
  LPM_q_ivl_36219 <= tmp_ivl_36221 & tmp_ivl_36217;
  new_AGEMA_signal_3025 <= tmp_ivl_36225(1);
  tmp_ivl_36223 <= tmp_ivl_36225(0);
  tmp_ivl_36225 <= LPM_d0_ivl_36229(0 + 1 downto 0);
  tmp_ivl_36230 <= new_AGEMA_signal_2790 & n3254;
  LPM_q_ivl_36233 <= tmp_ivl_36235 & tmp_ivl_36230;
  tmp_ivl_36237 <= new_AGEMA_signal_2859 & SboxInst_n345;
  LPM_q_ivl_36240 <= tmp_ivl_36242 & tmp_ivl_36237;
  tmp_ivl_36245 <= fresh(39);
  LPM_q_ivl_36247 <= tmp_ivl_36249 & tmp_ivl_36245;
  new_AGEMA_signal_3026 <= tmp_ivl_36253(1);
  tmp_ivl_36251 <= tmp_ivl_36253(0);
  tmp_ivl_36253 <= LPM_d0_ivl_36257(0 + 1 downto 0);
  tmp_ivl_36258 <= new_AGEMA_signal_2793 & n3253;
  LPM_q_ivl_36261 <= tmp_ivl_36263 & tmp_ivl_36258;
  tmp_ivl_36265 <= new_AGEMA_signal_2877 & SboxInst_n344;
  LPM_q_ivl_36268 <= tmp_ivl_36270 & tmp_ivl_36265;
  tmp_ivl_36273 <= fresh(40);
  LPM_q_ivl_36275 <= tmp_ivl_36277 & tmp_ivl_36273;
  new_AGEMA_signal_3027 <= tmp_ivl_36281(1);
  tmp_ivl_36279 <= tmp_ivl_36281(0);
  tmp_ivl_36281 <= LPM_d0_ivl_36285(0 + 1 downto 0);
  tmp_ivl_36286 <= new_AGEMA_signal_2795 & n3252;
  LPM_q_ivl_36289 <= tmp_ivl_36291 & tmp_ivl_36286;
  tmp_ivl_36293 <= new_AGEMA_signal_2875 & SboxInst_n343;
  LPM_q_ivl_36296 <= tmp_ivl_36298 & tmp_ivl_36293;
  tmp_ivl_36301 <= fresh(41);
  LPM_q_ivl_36303 <= tmp_ivl_36305 & tmp_ivl_36301;
  new_AGEMA_signal_3028 <= tmp_ivl_36309(1);
  tmp_ivl_36307 <= tmp_ivl_36309(0);
  tmp_ivl_36309 <= LPM_d0_ivl_36313(0 + 1 downto 0);
  tmp_ivl_36314 <= new_AGEMA_signal_2797 & n3251;
  LPM_q_ivl_36317 <= tmp_ivl_36319 & tmp_ivl_36314;
  tmp_ivl_36321 <= new_AGEMA_signal_2873 & SboxInst_n342;
  LPM_q_ivl_36324 <= tmp_ivl_36326 & tmp_ivl_36321;
  tmp_ivl_36329 <= fresh(42);
  LPM_q_ivl_36331 <= tmp_ivl_36333 & tmp_ivl_36329;
  new_AGEMA_signal_3029 <= tmp_ivl_36337(1);
  tmp_ivl_36335 <= tmp_ivl_36337(0);
  tmp_ivl_36337 <= LPM_d0_ivl_36341(0 + 1 downto 0);
  tmp_ivl_36342 <= new_AGEMA_signal_2800 & n3250;
  LPM_q_ivl_36345 <= tmp_ivl_36347 & tmp_ivl_36342;
  tmp_ivl_36349 <= new_AGEMA_signal_2880 & SboxInst_n341;
  LPM_q_ivl_36352 <= tmp_ivl_36354 & tmp_ivl_36349;
  tmp_ivl_36357 <= fresh(43);
  LPM_q_ivl_36359 <= tmp_ivl_36361 & tmp_ivl_36357;
  new_AGEMA_signal_3030 <= tmp_ivl_36365(1);
  tmp_ivl_36363 <= tmp_ivl_36365(0);
  tmp_ivl_36365 <= LPM_d0_ivl_36369(0 + 1 downto 0);
  tmp_ivl_36370 <= new_AGEMA_signal_2990 & n3232;
  LPM_q_ivl_36373 <= tmp_ivl_36375 & tmp_ivl_36370;
  tmp_ivl_36377 <= new_AGEMA_signal_2892 & SboxInst_n340;
  LPM_q_ivl_36380 <= tmp_ivl_36382 & tmp_ivl_36377;
  tmp_ivl_36385 <= fresh(44);
  LPM_q_ivl_36387 <= tmp_ivl_36389 & tmp_ivl_36385;
  new_AGEMA_signal_3518 <= tmp_ivl_36393(1);
  tmp_ivl_36391 <= tmp_ivl_36393(0);
  tmp_ivl_36393 <= LPM_d0_ivl_36397(0 + 1 downto 0);
  tmp_ivl_36398 <= new_AGEMA_signal_2803 & n3249;
  LPM_q_ivl_36401 <= tmp_ivl_36403 & tmp_ivl_36398;
  tmp_ivl_36405 <= new_AGEMA_signal_2879 & SboxInst_n339;
  LPM_q_ivl_36408 <= tmp_ivl_36410 & tmp_ivl_36405;
  tmp_ivl_36413 <= fresh(45);
  LPM_q_ivl_36415 <= tmp_ivl_36417 & tmp_ivl_36413;
  new_AGEMA_signal_3031 <= tmp_ivl_36421(1);
  tmp_ivl_36419 <= tmp_ivl_36421(0);
  tmp_ivl_36421 <= LPM_d0_ivl_36425(0 + 1 downto 0);
  tmp_ivl_36426 <= new_AGEMA_signal_2805 & n3248;
  LPM_q_ivl_36429 <= tmp_ivl_36431 & tmp_ivl_36426;
  tmp_ivl_36433 <= new_AGEMA_signal_2878 & SboxInst_n338;
  LPM_q_ivl_36436 <= tmp_ivl_36438 & tmp_ivl_36433;
  tmp_ivl_36441 <= fresh(46);
  LPM_q_ivl_36443 <= tmp_ivl_36445 & tmp_ivl_36441;
  new_AGEMA_signal_3032 <= tmp_ivl_36449(1);
  tmp_ivl_36447 <= tmp_ivl_36449(0);
  tmp_ivl_36449 <= LPM_d0_ivl_36453(0 + 1 downto 0);
  tmp_ivl_36454 <= new_AGEMA_signal_2807 & n3247;
  LPM_q_ivl_36457 <= tmp_ivl_36459 & tmp_ivl_36454;
  tmp_ivl_36461 <= new_AGEMA_signal_2876 & SboxInst_n337;
  LPM_q_ivl_36464 <= tmp_ivl_36466 & tmp_ivl_36461;
  tmp_ivl_36469 <= fresh(47);
  LPM_q_ivl_36471 <= tmp_ivl_36473 & tmp_ivl_36469;
  new_AGEMA_signal_3033 <= tmp_ivl_36477(1);
  tmp_ivl_36475 <= tmp_ivl_36477(0);
  tmp_ivl_36477 <= LPM_d0_ivl_36481(0 + 1 downto 0);
  tmp_ivl_36482 <= new_AGEMA_signal_2810 & n3246;
  LPM_q_ivl_36485 <= tmp_ivl_36487 & tmp_ivl_36482;
  tmp_ivl_36489 <= new_AGEMA_signal_2874 & SboxInst_n336;
  LPM_q_ivl_36492 <= tmp_ivl_36494 & tmp_ivl_36489;
  tmp_ivl_36497 <= fresh(48);
  LPM_q_ivl_36499 <= tmp_ivl_36501 & tmp_ivl_36497;
  new_AGEMA_signal_3034 <= tmp_ivl_36505(1);
  tmp_ivl_36503 <= tmp_ivl_36505(0);
  tmp_ivl_36505 <= LPM_d0_ivl_36509(0 + 1 downto 0);
  tmp_ivl_36510 <= new_AGEMA_signal_2813 & n3245;
  LPM_q_ivl_36513 <= tmp_ivl_36515 & tmp_ivl_36510;
  tmp_ivl_36517 <= new_AGEMA_signal_2884 & SboxInst_n335;
  LPM_q_ivl_36520 <= tmp_ivl_36522 & tmp_ivl_36517;
  tmp_ivl_36525 <= fresh(49);
  LPM_q_ivl_36527 <= tmp_ivl_36529 & tmp_ivl_36525;
  new_AGEMA_signal_3035 <= tmp_ivl_36533(1);
  tmp_ivl_36531 <= tmp_ivl_36533(0);
  tmp_ivl_36533 <= LPM_d0_ivl_36537(0 + 1 downto 0);
  tmp_ivl_36538 <= new_AGEMA_signal_2816 & n3244;
  LPM_q_ivl_36541 <= tmp_ivl_36543 & tmp_ivl_36538;
  tmp_ivl_36545 <= new_AGEMA_signal_2881 & SboxInst_n334;
  LPM_q_ivl_36548 <= tmp_ivl_36550 & tmp_ivl_36545;
  tmp_ivl_36553 <= fresh(50);
  LPM_q_ivl_36555 <= tmp_ivl_36557 & tmp_ivl_36553;
  new_AGEMA_signal_3036 <= tmp_ivl_36561(1);
  tmp_ivl_36559 <= tmp_ivl_36561(0);
  tmp_ivl_36561 <= LPM_d0_ivl_36565(0 + 1 downto 0);
  tmp_ivl_36566 <= new_AGEMA_signal_2819 & n3243;
  LPM_q_ivl_36569 <= tmp_ivl_36571 & tmp_ivl_36566;
  tmp_ivl_36573 <= new_AGEMA_signal_2883 & SboxInst_n333;
  LPM_q_ivl_36576 <= tmp_ivl_36578 & tmp_ivl_36573;
  tmp_ivl_36581 <= fresh(51);
  LPM_q_ivl_36583 <= tmp_ivl_36585 & tmp_ivl_36581;
  new_AGEMA_signal_3037 <= tmp_ivl_36589(1);
  tmp_ivl_36587 <= tmp_ivl_36589(0);
  tmp_ivl_36589 <= LPM_d0_ivl_36593(0 + 1 downto 0);
  tmp_ivl_36594 <= new_AGEMA_signal_2821 & n3242;
  LPM_q_ivl_36597 <= tmp_ivl_36599 & tmp_ivl_36594;
  tmp_ivl_36601 <= new_AGEMA_signal_2888 & SboxInst_n332;
  LPM_q_ivl_36604 <= tmp_ivl_36606 & tmp_ivl_36601;
  tmp_ivl_36609 <= fresh(52);
  LPM_q_ivl_36611 <= tmp_ivl_36613 & tmp_ivl_36609;
  new_AGEMA_signal_3038 <= tmp_ivl_36617(1);
  tmp_ivl_36615 <= tmp_ivl_36617(0);
  tmp_ivl_36617 <= LPM_d0_ivl_36621(0 + 1 downto 0);
  tmp_ivl_36622 <= new_AGEMA_signal_2823 & n3241;
  LPM_q_ivl_36625 <= tmp_ivl_36627 & tmp_ivl_36622;
  tmp_ivl_36629 <= new_AGEMA_signal_2887 & SboxInst_n331;
  LPM_q_ivl_36632 <= tmp_ivl_36634 & tmp_ivl_36629;
  tmp_ivl_36637 <= fresh(53);
  LPM_q_ivl_36639 <= tmp_ivl_36641 & tmp_ivl_36637;
  new_AGEMA_signal_3039 <= tmp_ivl_36645(1);
  tmp_ivl_36643 <= tmp_ivl_36645(0);
  tmp_ivl_36645 <= LPM_d0_ivl_36649(0 + 1 downto 0);
  tmp_ivl_36650 <= new_AGEMA_signal_2825 & n3240;
  LPM_q_ivl_36653 <= tmp_ivl_36655 & tmp_ivl_36650;
  tmp_ivl_36657 <= new_AGEMA_signal_2886 & SboxInst_n330;
  LPM_q_ivl_36660 <= tmp_ivl_36662 & tmp_ivl_36657;
  tmp_ivl_36665 <= fresh(54);
  LPM_q_ivl_36667 <= tmp_ivl_36669 & tmp_ivl_36665;
  new_AGEMA_signal_3040 <= tmp_ivl_36673(1);
  tmp_ivl_36671 <= tmp_ivl_36673(0);
  tmp_ivl_36673 <= LPM_d0_ivl_36677(0 + 1 downto 0);
  tmp_ivl_36678 <= new_AGEMA_signal_3515 & n3231;
  LPM_q_ivl_36681 <= tmp_ivl_36683 & tmp_ivl_36678;
  tmp_ivl_36685 <= new_AGEMA_signal_2891 & SboxInst_n329;
  LPM_q_ivl_36688 <= tmp_ivl_36690 & tmp_ivl_36685;
  tmp_ivl_36693 <= fresh(55);
  LPM_q_ivl_36695 <= tmp_ivl_36697 & tmp_ivl_36693;
  new_AGEMA_signal_3888 <= tmp_ivl_36701(1);
  tmp_ivl_36699 <= tmp_ivl_36701(0);
  tmp_ivl_36701 <= LPM_d0_ivl_36705(0 + 1 downto 0);
  tmp_ivl_36706 <= new_AGEMA_signal_2828 & n3238;
  LPM_q_ivl_36709 <= tmp_ivl_36711 & tmp_ivl_36706;
  tmp_ivl_36713 <= new_AGEMA_signal_2885 & SboxInst_n328;
  LPM_q_ivl_36716 <= tmp_ivl_36718 & tmp_ivl_36713;
  tmp_ivl_36721 <= fresh(56);
  LPM_q_ivl_36723 <= tmp_ivl_36725 & tmp_ivl_36721;
  new_AGEMA_signal_3041 <= tmp_ivl_36729(1);
  tmp_ivl_36727 <= tmp_ivl_36729(0);
  tmp_ivl_36729 <= LPM_d0_ivl_36733(0 + 1 downto 0);
  tmp_ivl_36734 <= new_AGEMA_signal_2837 & n3236;
  LPM_q_ivl_36737 <= tmp_ivl_36739 & tmp_ivl_36734;
  tmp_ivl_36741 <= new_AGEMA_signal_2882 & SboxInst_n327;
  LPM_q_ivl_36744 <= tmp_ivl_36746 & tmp_ivl_36741;
  tmp_ivl_36749 <= fresh(57);
  LPM_q_ivl_36751 <= tmp_ivl_36753 & tmp_ivl_36749;
  new_AGEMA_signal_3042 <= tmp_ivl_36757(1);
  tmp_ivl_36755 <= tmp_ivl_36757(0);
  tmp_ivl_36757 <= LPM_d0_ivl_36761(0 + 1 downto 0);
  tmp_ivl_36762 <= new_AGEMA_signal_2840 & n3235;
  LPM_q_ivl_36765 <= tmp_ivl_36767 & tmp_ivl_36762;
  tmp_ivl_36769 <= new_AGEMA_signal_2893 & SboxInst_n326;
  LPM_q_ivl_36772 <= tmp_ivl_36774 & tmp_ivl_36769;
  tmp_ivl_36777 <= fresh(58);
  LPM_q_ivl_36779 <= tmp_ivl_36781 & tmp_ivl_36777;
  new_AGEMA_signal_3043 <= tmp_ivl_36785(1);
  tmp_ivl_36783 <= tmp_ivl_36785(0);
  tmp_ivl_36785 <= LPM_d0_ivl_36789(0 + 1 downto 0);
  tmp_ivl_36790 <= new_AGEMA_signal_2846 & n3234;
  LPM_q_ivl_36793 <= tmp_ivl_36795 & tmp_ivl_36790;
  tmp_ivl_36797 <= new_AGEMA_signal_2889 & SboxInst_n325;
  LPM_q_ivl_36800 <= tmp_ivl_36802 & tmp_ivl_36797;
  tmp_ivl_36805 <= fresh(59);
  LPM_q_ivl_36807 <= tmp_ivl_36809 & tmp_ivl_36805;
  new_AGEMA_signal_3044 <= tmp_ivl_36813(1);
  tmp_ivl_36811 <= tmp_ivl_36813(0);
  tmp_ivl_36813 <= LPM_d0_ivl_36817(0 + 1 downto 0);
  tmp_ivl_36818 <= new_AGEMA_signal_3826 & n3230;
  LPM_q_ivl_36821 <= tmp_ivl_36823 & tmp_ivl_36818;
  tmp_ivl_36825 <= new_AGEMA_signal_2966 & SboxInst_n324;
  LPM_q_ivl_36828 <= tmp_ivl_36830 & tmp_ivl_36825;
  tmp_ivl_36833 <= fresh(60);
  LPM_q_ivl_36835 <= tmp_ivl_36837 & tmp_ivl_36833;
  new_AGEMA_signal_4201 <= tmp_ivl_36841(1);
  tmp_ivl_36839 <= tmp_ivl_36841(0);
  tmp_ivl_36841 <= LPM_d0_ivl_36845(0 + 1 downto 0);
  tmp_ivl_36846 <= new_AGEMA_signal_4433 & n3239;
  LPM_q_ivl_36849 <= tmp_ivl_36851 & tmp_ivl_36846;
  tmp_ivl_36853 <= new_AGEMA_signal_2963 & SboxInst_n323;
  LPM_q_ivl_36856 <= tmp_ivl_36858 & tmp_ivl_36853;
  tmp_ivl_36861 <= fresh(61);
  LPM_q_ivl_36863 <= tmp_ivl_36865 & tmp_ivl_36861;
  new_AGEMA_signal_4578 <= tmp_ivl_36869(1);
  tmp_ivl_36867 <= tmp_ivl_36869(0);
  tmp_ivl_36869 <= LPM_d0_ivl_36873(0 + 1 downto 0);
  tmp_ivl_36874 <= new_AGEMA_signal_2834 & n3237;
  LPM_q_ivl_36877 <= tmp_ivl_36879 & tmp_ivl_36874;
  tmp_ivl_36881 <= new_AGEMA_signal_2988 & SboxInst_n322;
  LPM_q_ivl_36884 <= tmp_ivl_36886 & tmp_ivl_36881;
  tmp_ivl_36889 <= fresh(62);
  LPM_q_ivl_36891 <= tmp_ivl_36893 & tmp_ivl_36889;
  new_AGEMA_signal_3045 <= tmp_ivl_36897(1);
  tmp_ivl_36895 <= tmp_ivl_36897(0);
  tmp_ivl_36897 <= LPM_d0_ivl_36901(0 + 1 downto 0);
  tmp_ivl_36902 <= new_AGEMA_signal_2692 & n3291;
  LPM_q_ivl_36905 <= tmp_ivl_36907 & tmp_ivl_36902;
  tmp_ivl_36909 <= new_AGEMA_signal_2986 & SboxInst_n321;
  LPM_q_ivl_36912 <= tmp_ivl_36914 & tmp_ivl_36909;
  tmp_ivl_36917 <= fresh(63);
  LPM_q_ivl_36919 <= tmp_ivl_36921 & tmp_ivl_36917;
  new_AGEMA_signal_3046 <= tmp_ivl_36925(1);
  tmp_ivl_36923 <= tmp_ivl_36925(0);
  tmp_ivl_36925 <= LPM_d0_ivl_36929(0 + 1 downto 0);
  tmp_ivl_36931 <= y4(0);
  tmp_ivl_36932 <= new_AGEMA_signal_2527 & tmp_ivl_36931;
  LPM_q_ivl_36935 <= tmp_ivl_36937 & tmp_ivl_36932;
  tmp_ivl_36939 <= new_AGEMA_signal_3047 & SboxInst_n320;
  LPM_q_ivl_36942 <= tmp_ivl_36944 & tmp_ivl_36939;
  tmp_ivl_36947 <= fresh(64);
  LPM_q_ivl_36949 <= tmp_ivl_36951 & tmp_ivl_36947;
  new_AGEMA_signal_3519 <= tmp_ivl_36955(1);
  tmp_ivl_36953 <= tmp_ivl_36955(0);
  tmp_ivl_36955 <= LPM_d0_ivl_36959(0 + 1 downto 0);
  tmp_ivl_36961 <= y4(10);
  tmp_ivl_36962 <= new_AGEMA_signal_2524 & tmp_ivl_36961;
  LPM_q_ivl_36965 <= tmp_ivl_36967 & tmp_ivl_36962;
  tmp_ivl_36969 <= new_AGEMA_signal_3048 & SboxInst_n319;
  LPM_q_ivl_36972 <= tmp_ivl_36974 & tmp_ivl_36969;
  tmp_ivl_36977 <= fresh(65);
  LPM_q_ivl_36979 <= tmp_ivl_36981 & tmp_ivl_36977;
  new_AGEMA_signal_3520 <= tmp_ivl_36985(1);
  tmp_ivl_36983 <= tmp_ivl_36985(0);
  tmp_ivl_36985 <= LPM_d0_ivl_36989(0 + 1 downto 0);
  tmp_ivl_36991 <= y4(11);
  tmp_ivl_36992 <= new_AGEMA_signal_2521 & tmp_ivl_36991;
  LPM_q_ivl_36995 <= tmp_ivl_36997 & tmp_ivl_36992;
  tmp_ivl_36999 <= new_AGEMA_signal_3049 & SboxInst_n318;
  LPM_q_ivl_37002 <= tmp_ivl_37004 & tmp_ivl_36999;
  tmp_ivl_37007 <= fresh(66);
  LPM_q_ivl_37009 <= tmp_ivl_37011 & tmp_ivl_37007;
  new_AGEMA_signal_3521 <= tmp_ivl_37015(1);
  tmp_ivl_37013 <= tmp_ivl_37015(0);
  tmp_ivl_37015 <= LPM_d0_ivl_37019(0 + 1 downto 0);
  tmp_ivl_37021 <= y4(12);
  tmp_ivl_37022 <= new_AGEMA_signal_2518 & tmp_ivl_37021;
  LPM_q_ivl_37025 <= tmp_ivl_37027 & tmp_ivl_37022;
  tmp_ivl_37029 <= new_AGEMA_signal_3050 & SboxInst_n317;
  LPM_q_ivl_37032 <= tmp_ivl_37034 & tmp_ivl_37029;
  tmp_ivl_37037 <= fresh(67);
  LPM_q_ivl_37039 <= tmp_ivl_37041 & tmp_ivl_37037;
  new_AGEMA_signal_3522 <= tmp_ivl_37045(1);
  tmp_ivl_37043 <= tmp_ivl_37045(0);
  tmp_ivl_37045 <= LPM_d0_ivl_37049(0 + 1 downto 0);
  tmp_ivl_37051 <= y4(13);
  tmp_ivl_37052 <= new_AGEMA_signal_2515 & tmp_ivl_37051;
  LPM_q_ivl_37055 <= tmp_ivl_37057 & tmp_ivl_37052;
  tmp_ivl_37059 <= new_AGEMA_signal_3051 & SboxInst_n316;
  LPM_q_ivl_37062 <= tmp_ivl_37064 & tmp_ivl_37059;
  tmp_ivl_37067 <= fresh(68);
  LPM_q_ivl_37069 <= tmp_ivl_37071 & tmp_ivl_37067;
  new_AGEMA_signal_3523 <= tmp_ivl_37075(1);
  tmp_ivl_37073 <= tmp_ivl_37075(0);
  tmp_ivl_37075 <= LPM_d0_ivl_37079(0 + 1 downto 0);
  tmp_ivl_37081 <= y4(14);
  tmp_ivl_37082 <= new_AGEMA_signal_2512 & tmp_ivl_37081;
  LPM_q_ivl_37085 <= tmp_ivl_37087 & tmp_ivl_37082;
  tmp_ivl_37089 <= new_AGEMA_signal_3052 & SboxInst_n315;
  LPM_q_ivl_37092 <= tmp_ivl_37094 & tmp_ivl_37089;
  tmp_ivl_37097 <= fresh(69);
  LPM_q_ivl_37099 <= tmp_ivl_37101 & tmp_ivl_37097;
  new_AGEMA_signal_3524 <= tmp_ivl_37105(1);
  tmp_ivl_37103 <= tmp_ivl_37105(0);
  tmp_ivl_37105 <= LPM_d0_ivl_37109(0 + 1 downto 0);
  tmp_ivl_37111 <= y4(15);
  tmp_ivl_37112 <= new_AGEMA_signal_2509 & tmp_ivl_37111;
  LPM_q_ivl_37115 <= tmp_ivl_37117 & tmp_ivl_37112;
  tmp_ivl_37119 <= new_AGEMA_signal_3053 & SboxInst_n314;
  LPM_q_ivl_37122 <= tmp_ivl_37124 & tmp_ivl_37119;
  tmp_ivl_37127 <= fresh(70);
  LPM_q_ivl_37129 <= tmp_ivl_37131 & tmp_ivl_37127;
  new_AGEMA_signal_3525 <= tmp_ivl_37135(1);
  tmp_ivl_37133 <= tmp_ivl_37135(0);
  tmp_ivl_37135 <= LPM_d0_ivl_37139(0 + 1 downto 0);
  tmp_ivl_37141 <= y4(16);
  tmp_ivl_37142 <= new_AGEMA_signal_2506 & tmp_ivl_37141;
  LPM_q_ivl_37145 <= tmp_ivl_37147 & tmp_ivl_37142;
  tmp_ivl_37149 <= new_AGEMA_signal_3054 & SboxInst_n313;
  LPM_q_ivl_37152 <= tmp_ivl_37154 & tmp_ivl_37149;
  tmp_ivl_37157 <= fresh(71);
  LPM_q_ivl_37159 <= tmp_ivl_37161 & tmp_ivl_37157;
  new_AGEMA_signal_3526 <= tmp_ivl_37165(1);
  tmp_ivl_37163 <= tmp_ivl_37165(0);
  tmp_ivl_37165 <= LPM_d0_ivl_37169(0 + 1 downto 0);
  tmp_ivl_37171 <= y4(17);
  tmp_ivl_37172 <= new_AGEMA_signal_2503 & tmp_ivl_37171;
  LPM_q_ivl_37175 <= tmp_ivl_37177 & tmp_ivl_37172;
  tmp_ivl_37179 <= new_AGEMA_signal_3055 & SboxInst_n312;
  LPM_q_ivl_37182 <= tmp_ivl_37184 & tmp_ivl_37179;
  tmp_ivl_37187 <= fresh(72);
  LPM_q_ivl_37189 <= tmp_ivl_37191 & tmp_ivl_37187;
  new_AGEMA_signal_3527 <= tmp_ivl_37195(1);
  tmp_ivl_37193 <= tmp_ivl_37195(0);
  tmp_ivl_37195 <= LPM_d0_ivl_37199(0 + 1 downto 0);
  tmp_ivl_37201 <= y4(18);
  tmp_ivl_37202 <= new_AGEMA_signal_2500 & tmp_ivl_37201;
  LPM_q_ivl_37205 <= tmp_ivl_37207 & tmp_ivl_37202;
  tmp_ivl_37209 <= new_AGEMA_signal_3056 & SboxInst_n311;
  LPM_q_ivl_37212 <= tmp_ivl_37214 & tmp_ivl_37209;
  tmp_ivl_37217 <= fresh(73);
  LPM_q_ivl_37219 <= tmp_ivl_37221 & tmp_ivl_37217;
  new_AGEMA_signal_3528 <= tmp_ivl_37225(1);
  tmp_ivl_37223 <= tmp_ivl_37225(0);
  tmp_ivl_37225 <= LPM_d0_ivl_37229(0 + 1 downto 0);
  tmp_ivl_37231 <= y4(19);
  tmp_ivl_37232 <= new_AGEMA_signal_2497 & tmp_ivl_37231;
  LPM_q_ivl_37235 <= tmp_ivl_37237 & tmp_ivl_37232;
  tmp_ivl_37239 <= new_AGEMA_signal_3057 & SboxInst_n310;
  LPM_q_ivl_37242 <= tmp_ivl_37244 & tmp_ivl_37239;
  tmp_ivl_37247 <= fresh(74);
  LPM_q_ivl_37249 <= tmp_ivl_37251 & tmp_ivl_37247;
  new_AGEMA_signal_3529 <= tmp_ivl_37255(1);
  tmp_ivl_37253 <= tmp_ivl_37255(0);
  tmp_ivl_37255 <= LPM_d0_ivl_37259(0 + 1 downto 0);
  tmp_ivl_37261 <= y4(1);
  tmp_ivl_37262 <= new_AGEMA_signal_2494 & tmp_ivl_37261;
  LPM_q_ivl_37265 <= tmp_ivl_37267 & tmp_ivl_37262;
  tmp_ivl_37269 <= new_AGEMA_signal_3058 & SboxInst_n309;
  LPM_q_ivl_37272 <= tmp_ivl_37274 & tmp_ivl_37269;
  tmp_ivl_37277 <= fresh(75);
  LPM_q_ivl_37279 <= tmp_ivl_37281 & tmp_ivl_37277;
  new_AGEMA_signal_3530 <= tmp_ivl_37285(1);
  tmp_ivl_37283 <= tmp_ivl_37285(0);
  tmp_ivl_37285 <= LPM_d0_ivl_37289(0 + 1 downto 0);
  tmp_ivl_37291 <= y4(20);
  tmp_ivl_37292 <= new_AGEMA_signal_2491 & tmp_ivl_37291;
  LPM_q_ivl_37295 <= tmp_ivl_37297 & tmp_ivl_37292;
  tmp_ivl_37299 <= new_AGEMA_signal_3059 & SboxInst_n308;
  LPM_q_ivl_37302 <= tmp_ivl_37304 & tmp_ivl_37299;
  tmp_ivl_37307 <= fresh(76);
  LPM_q_ivl_37309 <= tmp_ivl_37311 & tmp_ivl_37307;
  new_AGEMA_signal_3531 <= tmp_ivl_37315(1);
  tmp_ivl_37313 <= tmp_ivl_37315(0);
  tmp_ivl_37315 <= LPM_d0_ivl_37319(0 + 1 downto 0);
  tmp_ivl_37321 <= y4(21);
  tmp_ivl_37322 <= new_AGEMA_signal_2488 & tmp_ivl_37321;
  LPM_q_ivl_37325 <= tmp_ivl_37327 & tmp_ivl_37322;
  tmp_ivl_37329 <= new_AGEMA_signal_3060 & SboxInst_n307;
  LPM_q_ivl_37332 <= tmp_ivl_37334 & tmp_ivl_37329;
  tmp_ivl_37337 <= fresh(77);
  LPM_q_ivl_37339 <= tmp_ivl_37341 & tmp_ivl_37337;
  new_AGEMA_signal_3532 <= tmp_ivl_37345(1);
  tmp_ivl_37343 <= tmp_ivl_37345(0);
  tmp_ivl_37345 <= LPM_d0_ivl_37349(0 + 1 downto 0);
  tmp_ivl_37351 <= y4(22);
  tmp_ivl_37352 <= new_AGEMA_signal_2485 & tmp_ivl_37351;
  LPM_q_ivl_37355 <= tmp_ivl_37357 & tmp_ivl_37352;
  tmp_ivl_37359 <= new_AGEMA_signal_3061 & SboxInst_n306;
  LPM_q_ivl_37362 <= tmp_ivl_37364 & tmp_ivl_37359;
  tmp_ivl_37367 <= fresh(78);
  LPM_q_ivl_37369 <= tmp_ivl_37371 & tmp_ivl_37367;
  new_AGEMA_signal_3533 <= tmp_ivl_37375(1);
  tmp_ivl_37373 <= tmp_ivl_37375(0);
  tmp_ivl_37375 <= LPM_d0_ivl_37379(0 + 1 downto 0);
  tmp_ivl_37381 <= y4(23);
  tmp_ivl_37382 <= new_AGEMA_signal_2482 & tmp_ivl_37381;
  LPM_q_ivl_37385 <= tmp_ivl_37387 & tmp_ivl_37382;
  tmp_ivl_37389 <= new_AGEMA_signal_3062 & SboxInst_n305;
  LPM_q_ivl_37392 <= tmp_ivl_37394 & tmp_ivl_37389;
  tmp_ivl_37397 <= fresh(79);
  LPM_q_ivl_37399 <= tmp_ivl_37401 & tmp_ivl_37397;
  new_AGEMA_signal_3534 <= tmp_ivl_37405(1);
  tmp_ivl_37403 <= tmp_ivl_37405(0);
  tmp_ivl_37405 <= LPM_d0_ivl_37409(0 + 1 downto 0);
  tmp_ivl_37411 <= y4(24);
  tmp_ivl_37412 <= new_AGEMA_signal_2479 & tmp_ivl_37411;
  LPM_q_ivl_37415 <= tmp_ivl_37417 & tmp_ivl_37412;
  tmp_ivl_37419 <= new_AGEMA_signal_3063 & SboxInst_n304;
  LPM_q_ivl_37422 <= tmp_ivl_37424 & tmp_ivl_37419;
  tmp_ivl_37427 <= fresh(80);
  LPM_q_ivl_37429 <= tmp_ivl_37431 & tmp_ivl_37427;
  new_AGEMA_signal_3535 <= tmp_ivl_37435(1);
  tmp_ivl_37433 <= tmp_ivl_37435(0);
  tmp_ivl_37435 <= LPM_d0_ivl_37439(0 + 1 downto 0);
  tmp_ivl_37441 <= y4(25);
  tmp_ivl_37442 <= new_AGEMA_signal_2476 & tmp_ivl_37441;
  LPM_q_ivl_37445 <= tmp_ivl_37447 & tmp_ivl_37442;
  tmp_ivl_37449 <= new_AGEMA_signal_3064 & SboxInst_n303;
  LPM_q_ivl_37452 <= tmp_ivl_37454 & tmp_ivl_37449;
  tmp_ivl_37457 <= fresh(81);
  LPM_q_ivl_37459 <= tmp_ivl_37461 & tmp_ivl_37457;
  new_AGEMA_signal_3536 <= tmp_ivl_37465(1);
  tmp_ivl_37463 <= tmp_ivl_37465(0);
  tmp_ivl_37465 <= LPM_d0_ivl_37469(0 + 1 downto 0);
  tmp_ivl_37471 <= y4(26);
  tmp_ivl_37472 <= new_AGEMA_signal_2473 & tmp_ivl_37471;
  LPM_q_ivl_37475 <= tmp_ivl_37477 & tmp_ivl_37472;
  tmp_ivl_37479 <= new_AGEMA_signal_3065 & SboxInst_n302;
  LPM_q_ivl_37482 <= tmp_ivl_37484 & tmp_ivl_37479;
  tmp_ivl_37487 <= fresh(82);
  LPM_q_ivl_37489 <= tmp_ivl_37491 & tmp_ivl_37487;
  new_AGEMA_signal_3537 <= tmp_ivl_37495(1);
  tmp_ivl_37493 <= tmp_ivl_37495(0);
  tmp_ivl_37495 <= LPM_d0_ivl_37499(0 + 1 downto 0);
  tmp_ivl_37501 <= y4(27);
  tmp_ivl_37502 <= new_AGEMA_signal_2470 & tmp_ivl_37501;
  LPM_q_ivl_37505 <= tmp_ivl_37507 & tmp_ivl_37502;
  tmp_ivl_37509 <= new_AGEMA_signal_3066 & SboxInst_n301;
  LPM_q_ivl_37512 <= tmp_ivl_37514 & tmp_ivl_37509;
  tmp_ivl_37517 <= fresh(83);
  LPM_q_ivl_37519 <= tmp_ivl_37521 & tmp_ivl_37517;
  new_AGEMA_signal_3538 <= tmp_ivl_37525(1);
  tmp_ivl_37523 <= tmp_ivl_37525(0);
  tmp_ivl_37525 <= LPM_d0_ivl_37529(0 + 1 downto 0);
  tmp_ivl_37531 <= y4(28);
  tmp_ivl_37532 <= new_AGEMA_signal_2467 & tmp_ivl_37531;
  LPM_q_ivl_37535 <= tmp_ivl_37537 & tmp_ivl_37532;
  tmp_ivl_37539 <= new_AGEMA_signal_3067 & SboxInst_n300;
  LPM_q_ivl_37542 <= tmp_ivl_37544 & tmp_ivl_37539;
  tmp_ivl_37547 <= fresh(84);
  LPM_q_ivl_37549 <= tmp_ivl_37551 & tmp_ivl_37547;
  new_AGEMA_signal_3539 <= tmp_ivl_37555(1);
  tmp_ivl_37553 <= tmp_ivl_37555(0);
  tmp_ivl_37555 <= LPM_d0_ivl_37559(0 + 1 downto 0);
  tmp_ivl_37561 <= y4(29);
  tmp_ivl_37562 <= new_AGEMA_signal_2464 & tmp_ivl_37561;
  LPM_q_ivl_37565 <= tmp_ivl_37567 & tmp_ivl_37562;
  tmp_ivl_37569 <= new_AGEMA_signal_3068 & SboxInst_n299;
  LPM_q_ivl_37572 <= tmp_ivl_37574 & tmp_ivl_37569;
  tmp_ivl_37577 <= fresh(85);
  LPM_q_ivl_37579 <= tmp_ivl_37581 & tmp_ivl_37577;
  new_AGEMA_signal_3540 <= tmp_ivl_37585(1);
  tmp_ivl_37583 <= tmp_ivl_37585(0);
  tmp_ivl_37585 <= LPM_d0_ivl_37589(0 + 1 downto 0);
  tmp_ivl_37591 <= y4(2);
  tmp_ivl_37592 <= new_AGEMA_signal_2461 & tmp_ivl_37591;
  LPM_q_ivl_37595 <= tmp_ivl_37597 & tmp_ivl_37592;
  tmp_ivl_37599 <= new_AGEMA_signal_3069 & SboxInst_n298;
  LPM_q_ivl_37602 <= tmp_ivl_37604 & tmp_ivl_37599;
  tmp_ivl_37607 <= fresh(86);
  LPM_q_ivl_37609 <= tmp_ivl_37611 & tmp_ivl_37607;
  new_AGEMA_signal_3541 <= tmp_ivl_37615(1);
  tmp_ivl_37613 <= tmp_ivl_37615(0);
  tmp_ivl_37615 <= LPM_d0_ivl_37619(0 + 1 downto 0);
  tmp_ivl_37621 <= y4(30);
  tmp_ivl_37622 <= new_AGEMA_signal_2458 & tmp_ivl_37621;
  LPM_q_ivl_37625 <= tmp_ivl_37627 & tmp_ivl_37622;
  tmp_ivl_37629 <= new_AGEMA_signal_3070 & SboxInst_n297;
  LPM_q_ivl_37632 <= tmp_ivl_37634 & tmp_ivl_37629;
  tmp_ivl_37637 <= fresh(87);
  LPM_q_ivl_37639 <= tmp_ivl_37641 & tmp_ivl_37637;
  new_AGEMA_signal_3542 <= tmp_ivl_37645(1);
  tmp_ivl_37643 <= tmp_ivl_37645(0);
  tmp_ivl_37645 <= LPM_d0_ivl_37649(0 + 1 downto 0);
  tmp_ivl_37651 <= y4(31);
  tmp_ivl_37652 <= new_AGEMA_signal_2455 & tmp_ivl_37651;
  LPM_q_ivl_37655 <= tmp_ivl_37657 & tmp_ivl_37652;
  tmp_ivl_37659 <= new_AGEMA_signal_3071 & SboxInst_n296;
  LPM_q_ivl_37662 <= tmp_ivl_37664 & tmp_ivl_37659;
  tmp_ivl_37667 <= fresh(88);
  LPM_q_ivl_37669 <= tmp_ivl_37671 & tmp_ivl_37667;
  new_AGEMA_signal_3543 <= tmp_ivl_37675(1);
  tmp_ivl_37673 <= tmp_ivl_37675(0);
  tmp_ivl_37675 <= LPM_d0_ivl_37679(0 + 1 downto 0);
  tmp_ivl_37681 <= y4(32);
  tmp_ivl_37682 <= new_AGEMA_signal_2452 & tmp_ivl_37681;
  LPM_q_ivl_37685 <= tmp_ivl_37687 & tmp_ivl_37682;
  tmp_ivl_37689 <= new_AGEMA_signal_3072 & SboxInst_n295;
  LPM_q_ivl_37692 <= tmp_ivl_37694 & tmp_ivl_37689;
  tmp_ivl_37697 <= fresh(89);
  LPM_q_ivl_37699 <= tmp_ivl_37701 & tmp_ivl_37697;
  new_AGEMA_signal_3544 <= tmp_ivl_37705(1);
  tmp_ivl_37703 <= tmp_ivl_37705(0);
  tmp_ivl_37705 <= LPM_d0_ivl_37709(0 + 1 downto 0);
  tmp_ivl_37711 <= y4(33);
  tmp_ivl_37712 <= new_AGEMA_signal_2449 & tmp_ivl_37711;
  LPM_q_ivl_37715 <= tmp_ivl_37717 & tmp_ivl_37712;
  tmp_ivl_37719 <= new_AGEMA_signal_3073 & SboxInst_n294;
  LPM_q_ivl_37722 <= tmp_ivl_37724 & tmp_ivl_37719;
  tmp_ivl_37727 <= fresh(90);
  LPM_q_ivl_37729 <= tmp_ivl_37731 & tmp_ivl_37727;
  new_AGEMA_signal_3545 <= tmp_ivl_37735(1);
  tmp_ivl_37733 <= tmp_ivl_37735(0);
  tmp_ivl_37735 <= LPM_d0_ivl_37739(0 + 1 downto 0);
  tmp_ivl_37741 <= y4(34);
  tmp_ivl_37742 <= new_AGEMA_signal_2446 & tmp_ivl_37741;
  LPM_q_ivl_37745 <= tmp_ivl_37747 & tmp_ivl_37742;
  tmp_ivl_37749 <= new_AGEMA_signal_3074 & SboxInst_n293;
  LPM_q_ivl_37752 <= tmp_ivl_37754 & tmp_ivl_37749;
  tmp_ivl_37757 <= fresh(91);
  LPM_q_ivl_37759 <= tmp_ivl_37761 & tmp_ivl_37757;
  new_AGEMA_signal_3546 <= tmp_ivl_37765(1);
  tmp_ivl_37763 <= tmp_ivl_37765(0);
  tmp_ivl_37765 <= LPM_d0_ivl_37769(0 + 1 downto 0);
  tmp_ivl_37771 <= y4(35);
  tmp_ivl_37772 <= new_AGEMA_signal_2443 & tmp_ivl_37771;
  LPM_q_ivl_37775 <= tmp_ivl_37777 & tmp_ivl_37772;
  tmp_ivl_37779 <= new_AGEMA_signal_3075 & SboxInst_n292;
  LPM_q_ivl_37782 <= tmp_ivl_37784 & tmp_ivl_37779;
  tmp_ivl_37787 <= fresh(92);
  LPM_q_ivl_37789 <= tmp_ivl_37791 & tmp_ivl_37787;
  new_AGEMA_signal_3547 <= tmp_ivl_37795(1);
  tmp_ivl_37793 <= tmp_ivl_37795(0);
  tmp_ivl_37795 <= LPM_d0_ivl_37799(0 + 1 downto 0);
  tmp_ivl_37801 <= y4(36);
  tmp_ivl_37802 <= new_AGEMA_signal_2440 & tmp_ivl_37801;
  LPM_q_ivl_37805 <= tmp_ivl_37807 & tmp_ivl_37802;
  tmp_ivl_37809 <= new_AGEMA_signal_3076 & SboxInst_n291;
  LPM_q_ivl_37812 <= tmp_ivl_37814 & tmp_ivl_37809;
  tmp_ivl_37817 <= fresh(93);
  LPM_q_ivl_37819 <= tmp_ivl_37821 & tmp_ivl_37817;
  new_AGEMA_signal_3548 <= tmp_ivl_37825(1);
  tmp_ivl_37823 <= tmp_ivl_37825(0);
  tmp_ivl_37825 <= LPM_d0_ivl_37829(0 + 1 downto 0);
  tmp_ivl_37831 <= y4(37);
  tmp_ivl_37832 <= new_AGEMA_signal_2437 & tmp_ivl_37831;
  LPM_q_ivl_37835 <= tmp_ivl_37837 & tmp_ivl_37832;
  tmp_ivl_37839 <= new_AGEMA_signal_3077 & SboxInst_n290;
  LPM_q_ivl_37842 <= tmp_ivl_37844 & tmp_ivl_37839;
  tmp_ivl_37847 <= fresh(94);
  LPM_q_ivl_37849 <= tmp_ivl_37851 & tmp_ivl_37847;
  new_AGEMA_signal_3549 <= tmp_ivl_37855(1);
  tmp_ivl_37853 <= tmp_ivl_37855(0);
  tmp_ivl_37855 <= LPM_d0_ivl_37859(0 + 1 downto 0);
  tmp_ivl_37861 <= y4(38);
  tmp_ivl_37862 <= new_AGEMA_signal_2434 & tmp_ivl_37861;
  LPM_q_ivl_37865 <= tmp_ivl_37867 & tmp_ivl_37862;
  tmp_ivl_37869 <= new_AGEMA_signal_3078 & SboxInst_n289;
  LPM_q_ivl_37872 <= tmp_ivl_37874 & tmp_ivl_37869;
  tmp_ivl_37877 <= fresh(95);
  LPM_q_ivl_37879 <= tmp_ivl_37881 & tmp_ivl_37877;
  new_AGEMA_signal_3550 <= tmp_ivl_37885(1);
  tmp_ivl_37883 <= tmp_ivl_37885(0);
  tmp_ivl_37885 <= LPM_d0_ivl_37889(0 + 1 downto 0);
  tmp_ivl_37891 <= y4(39);
  tmp_ivl_37892 <= new_AGEMA_signal_2431 & tmp_ivl_37891;
  LPM_q_ivl_37895 <= tmp_ivl_37897 & tmp_ivl_37892;
  tmp_ivl_37899 <= new_AGEMA_signal_3079 & SboxInst_n288;
  LPM_q_ivl_37902 <= tmp_ivl_37904 & tmp_ivl_37899;
  tmp_ivl_37907 <= fresh(96);
  LPM_q_ivl_37909 <= tmp_ivl_37911 & tmp_ivl_37907;
  new_AGEMA_signal_3551 <= tmp_ivl_37915(1);
  tmp_ivl_37913 <= tmp_ivl_37915(0);
  tmp_ivl_37915 <= LPM_d0_ivl_37919(0 + 1 downto 0);
  tmp_ivl_37921 <= y4(3);
  tmp_ivl_37922 <= new_AGEMA_signal_2428 & tmp_ivl_37921;
  LPM_q_ivl_37925 <= tmp_ivl_37927 & tmp_ivl_37922;
  tmp_ivl_37929 <= new_AGEMA_signal_3080 & SboxInst_n287;
  LPM_q_ivl_37932 <= tmp_ivl_37934 & tmp_ivl_37929;
  tmp_ivl_37937 <= fresh(97);
  LPM_q_ivl_37939 <= tmp_ivl_37941 & tmp_ivl_37937;
  new_AGEMA_signal_3552 <= tmp_ivl_37945(1);
  tmp_ivl_37943 <= tmp_ivl_37945(0);
  tmp_ivl_37945 <= LPM_d0_ivl_37949(0 + 1 downto 0);
  tmp_ivl_37951 <= y4(40);
  tmp_ivl_37952 <= new_AGEMA_signal_2425 & tmp_ivl_37951;
  LPM_q_ivl_37955 <= tmp_ivl_37957 & tmp_ivl_37952;
  tmp_ivl_37959 <= new_AGEMA_signal_3081 & SboxInst_n286;
  LPM_q_ivl_37962 <= tmp_ivl_37964 & tmp_ivl_37959;
  tmp_ivl_37967 <= fresh(98);
  LPM_q_ivl_37969 <= tmp_ivl_37971 & tmp_ivl_37967;
  new_AGEMA_signal_3553 <= tmp_ivl_37975(1);
  tmp_ivl_37973 <= tmp_ivl_37975(0);
  tmp_ivl_37975 <= LPM_d0_ivl_37979(0 + 1 downto 0);
  tmp_ivl_37981 <= y4(41);
  tmp_ivl_37982 <= new_AGEMA_signal_2422 & tmp_ivl_37981;
  LPM_q_ivl_37985 <= tmp_ivl_37987 & tmp_ivl_37982;
  tmp_ivl_37989 <= new_AGEMA_signal_3082 & SboxInst_n285;
  LPM_q_ivl_37992 <= tmp_ivl_37994 & tmp_ivl_37989;
  tmp_ivl_37997 <= fresh(99);
  LPM_q_ivl_37999 <= tmp_ivl_38001 & tmp_ivl_37997;
  new_AGEMA_signal_3554 <= tmp_ivl_38005(1);
  tmp_ivl_38003 <= tmp_ivl_38005(0);
  tmp_ivl_38005 <= LPM_d0_ivl_38009(0 + 1 downto 0);
  tmp_ivl_38011 <= y4(42);
  tmp_ivl_38012 <= new_AGEMA_signal_2419 & tmp_ivl_38011;
  LPM_q_ivl_38015 <= tmp_ivl_38017 & tmp_ivl_38012;
  tmp_ivl_38019 <= new_AGEMA_signal_3083 & SboxInst_n284;
  LPM_q_ivl_38022 <= tmp_ivl_38024 & tmp_ivl_38019;
  tmp_ivl_38027 <= fresh(100);
  LPM_q_ivl_38029 <= tmp_ivl_38031 & tmp_ivl_38027;
  new_AGEMA_signal_3555 <= tmp_ivl_38035(1);
  tmp_ivl_38033 <= tmp_ivl_38035(0);
  tmp_ivl_38035 <= LPM_d0_ivl_38039(0 + 1 downto 0);
  tmp_ivl_38041 <= y4(43);
  tmp_ivl_38042 <= new_AGEMA_signal_2416 & tmp_ivl_38041;
  LPM_q_ivl_38045 <= tmp_ivl_38047 & tmp_ivl_38042;
  tmp_ivl_38049 <= new_AGEMA_signal_3084 & SboxInst_n283;
  LPM_q_ivl_38052 <= tmp_ivl_38054 & tmp_ivl_38049;
  tmp_ivl_38057 <= fresh(101);
  LPM_q_ivl_38059 <= tmp_ivl_38061 & tmp_ivl_38057;
  new_AGEMA_signal_3556 <= tmp_ivl_38065(1);
  tmp_ivl_38063 <= tmp_ivl_38065(0);
  tmp_ivl_38065 <= LPM_d0_ivl_38069(0 + 1 downto 0);
  tmp_ivl_38071 <= y4(44);
  tmp_ivl_38072 <= new_AGEMA_signal_2413 & tmp_ivl_38071;
  LPM_q_ivl_38075 <= tmp_ivl_38077 & tmp_ivl_38072;
  tmp_ivl_38079 <= new_AGEMA_signal_3085 & SboxInst_n282;
  LPM_q_ivl_38082 <= tmp_ivl_38084 & tmp_ivl_38079;
  tmp_ivl_38087 <= fresh(102);
  LPM_q_ivl_38089 <= tmp_ivl_38091 & tmp_ivl_38087;
  new_AGEMA_signal_3557 <= tmp_ivl_38095(1);
  tmp_ivl_38093 <= tmp_ivl_38095(0);
  tmp_ivl_38095 <= LPM_d0_ivl_38099(0 + 1 downto 0);
  tmp_ivl_38101 <= y4(45);
  tmp_ivl_38102 <= new_AGEMA_signal_2410 & tmp_ivl_38101;
  LPM_q_ivl_38105 <= tmp_ivl_38107 & tmp_ivl_38102;
  tmp_ivl_38109 <= new_AGEMA_signal_3086 & SboxInst_n281;
  LPM_q_ivl_38112 <= tmp_ivl_38114 & tmp_ivl_38109;
  tmp_ivl_38117 <= fresh(103);
  LPM_q_ivl_38119 <= tmp_ivl_38121 & tmp_ivl_38117;
  new_AGEMA_signal_3558 <= tmp_ivl_38125(1);
  tmp_ivl_38123 <= tmp_ivl_38125(0);
  tmp_ivl_38125 <= LPM_d0_ivl_38129(0 + 1 downto 0);
  tmp_ivl_38131 <= y4(46);
  tmp_ivl_38132 <= new_AGEMA_signal_2407 & tmp_ivl_38131;
  LPM_q_ivl_38135 <= tmp_ivl_38137 & tmp_ivl_38132;
  tmp_ivl_38139 <= new_AGEMA_signal_3087 & SboxInst_n280;
  LPM_q_ivl_38142 <= tmp_ivl_38144 & tmp_ivl_38139;
  tmp_ivl_38147 <= fresh(104);
  LPM_q_ivl_38149 <= tmp_ivl_38151 & tmp_ivl_38147;
  new_AGEMA_signal_3559 <= tmp_ivl_38155(1);
  tmp_ivl_38153 <= tmp_ivl_38155(0);
  tmp_ivl_38155 <= LPM_d0_ivl_38159(0 + 1 downto 0);
  tmp_ivl_38161 <= y4(47);
  tmp_ivl_38162 <= new_AGEMA_signal_2404 & tmp_ivl_38161;
  LPM_q_ivl_38165 <= tmp_ivl_38167 & tmp_ivl_38162;
  tmp_ivl_38169 <= new_AGEMA_signal_3088 & SboxInst_n279;
  LPM_q_ivl_38172 <= tmp_ivl_38174 & tmp_ivl_38169;
  tmp_ivl_38177 <= fresh(105);
  LPM_q_ivl_38179 <= tmp_ivl_38181 & tmp_ivl_38177;
  new_AGEMA_signal_3560 <= tmp_ivl_38185(1);
  tmp_ivl_38183 <= tmp_ivl_38185(0);
  tmp_ivl_38185 <= LPM_d0_ivl_38189(0 + 1 downto 0);
  tmp_ivl_38191 <= y4(48);
  tmp_ivl_38192 <= new_AGEMA_signal_2401 & tmp_ivl_38191;
  LPM_q_ivl_38195 <= tmp_ivl_38197 & tmp_ivl_38192;
  tmp_ivl_38199 <= new_AGEMA_signal_3089 & SboxInst_n278;
  LPM_q_ivl_38202 <= tmp_ivl_38204 & tmp_ivl_38199;
  tmp_ivl_38207 <= fresh(106);
  LPM_q_ivl_38209 <= tmp_ivl_38211 & tmp_ivl_38207;
  new_AGEMA_signal_3561 <= tmp_ivl_38215(1);
  tmp_ivl_38213 <= tmp_ivl_38215(0);
  tmp_ivl_38215 <= LPM_d0_ivl_38219(0 + 1 downto 0);
  tmp_ivl_38221 <= y4(49);
  tmp_ivl_38222 <= new_AGEMA_signal_2398 & tmp_ivl_38221;
  LPM_q_ivl_38225 <= tmp_ivl_38227 & tmp_ivl_38222;
  tmp_ivl_38229 <= new_AGEMA_signal_3090 & SboxInst_n277;
  LPM_q_ivl_38232 <= tmp_ivl_38234 & tmp_ivl_38229;
  tmp_ivl_38237 <= fresh(107);
  LPM_q_ivl_38239 <= tmp_ivl_38241 & tmp_ivl_38237;
  new_AGEMA_signal_3562 <= tmp_ivl_38245(1);
  tmp_ivl_38243 <= tmp_ivl_38245(0);
  tmp_ivl_38245 <= LPM_d0_ivl_38249(0 + 1 downto 0);
  tmp_ivl_38251 <= y4(4);
  tmp_ivl_38252 <= new_AGEMA_signal_2395 & tmp_ivl_38251;
  LPM_q_ivl_38255 <= tmp_ivl_38257 & tmp_ivl_38252;
  tmp_ivl_38259 <= new_AGEMA_signal_3091 & SboxInst_n276;
  LPM_q_ivl_38262 <= tmp_ivl_38264 & tmp_ivl_38259;
  tmp_ivl_38267 <= fresh(108);
  LPM_q_ivl_38269 <= tmp_ivl_38271 & tmp_ivl_38267;
  new_AGEMA_signal_3563 <= tmp_ivl_38275(1);
  tmp_ivl_38273 <= tmp_ivl_38275(0);
  tmp_ivl_38275 <= LPM_d0_ivl_38279(0 + 1 downto 0);
  tmp_ivl_38281 <= y4(50);
  tmp_ivl_38282 <= new_AGEMA_signal_2392 & tmp_ivl_38281;
  LPM_q_ivl_38285 <= tmp_ivl_38287 & tmp_ivl_38282;
  tmp_ivl_38289 <= new_AGEMA_signal_3092 & SboxInst_n275;
  LPM_q_ivl_38292 <= tmp_ivl_38294 & tmp_ivl_38289;
  tmp_ivl_38297 <= fresh(109);
  LPM_q_ivl_38299 <= tmp_ivl_38301 & tmp_ivl_38297;
  new_AGEMA_signal_3564 <= tmp_ivl_38305(1);
  tmp_ivl_38303 <= tmp_ivl_38305(0);
  tmp_ivl_38305 <= LPM_d0_ivl_38309(0 + 1 downto 0);
  tmp_ivl_38311 <= y4(51);
  tmp_ivl_38312 <= new_AGEMA_signal_2389 & tmp_ivl_38311;
  LPM_q_ivl_38315 <= tmp_ivl_38317 & tmp_ivl_38312;
  tmp_ivl_38319 <= new_AGEMA_signal_3093 & SboxInst_n274;
  LPM_q_ivl_38322 <= tmp_ivl_38324 & tmp_ivl_38319;
  tmp_ivl_38327 <= fresh(110);
  LPM_q_ivl_38329 <= tmp_ivl_38331 & tmp_ivl_38327;
  new_AGEMA_signal_3565 <= tmp_ivl_38335(1);
  tmp_ivl_38333 <= tmp_ivl_38335(0);
  tmp_ivl_38335 <= LPM_d0_ivl_38339(0 + 1 downto 0);
  tmp_ivl_38341 <= y4(52);
  tmp_ivl_38342 <= new_AGEMA_signal_2386 & tmp_ivl_38341;
  LPM_q_ivl_38345 <= tmp_ivl_38347 & tmp_ivl_38342;
  tmp_ivl_38349 <= new_AGEMA_signal_3094 & SboxInst_n273;
  LPM_q_ivl_38352 <= tmp_ivl_38354 & tmp_ivl_38349;
  tmp_ivl_38357 <= fresh(111);
  LPM_q_ivl_38359 <= tmp_ivl_38361 & tmp_ivl_38357;
  new_AGEMA_signal_3566 <= tmp_ivl_38365(1);
  tmp_ivl_38363 <= tmp_ivl_38365(0);
  tmp_ivl_38365 <= LPM_d0_ivl_38369(0 + 1 downto 0);
  tmp_ivl_38371 <= y4(53);
  tmp_ivl_38372 <= new_AGEMA_signal_2383 & tmp_ivl_38371;
  LPM_q_ivl_38375 <= tmp_ivl_38377 & tmp_ivl_38372;
  tmp_ivl_38379 <= new_AGEMA_signal_3095 & SboxInst_n272;
  LPM_q_ivl_38382 <= tmp_ivl_38384 & tmp_ivl_38379;
  tmp_ivl_38387 <= fresh(112);
  LPM_q_ivl_38389 <= tmp_ivl_38391 & tmp_ivl_38387;
  new_AGEMA_signal_3567 <= tmp_ivl_38395(1);
  tmp_ivl_38393 <= tmp_ivl_38395(0);
  tmp_ivl_38395 <= LPM_d0_ivl_38399(0 + 1 downto 0);
  tmp_ivl_38401 <= y4(54);
  tmp_ivl_38402 <= new_AGEMA_signal_2380 & tmp_ivl_38401;
  LPM_q_ivl_38405 <= tmp_ivl_38407 & tmp_ivl_38402;
  tmp_ivl_38409 <= new_AGEMA_signal_3096 & SboxInst_n271;
  LPM_q_ivl_38412 <= tmp_ivl_38414 & tmp_ivl_38409;
  tmp_ivl_38417 <= fresh(113);
  LPM_q_ivl_38419 <= tmp_ivl_38421 & tmp_ivl_38417;
  new_AGEMA_signal_3568 <= tmp_ivl_38425(1);
  tmp_ivl_38423 <= tmp_ivl_38425(0);
  tmp_ivl_38425 <= LPM_d0_ivl_38429(0 + 1 downto 0);
  tmp_ivl_38431 <= y4(55);
  tmp_ivl_38432 <= new_AGEMA_signal_2377 & tmp_ivl_38431;
  LPM_q_ivl_38435 <= tmp_ivl_38437 & tmp_ivl_38432;
  tmp_ivl_38439 <= new_AGEMA_signal_3097 & SboxInst_n270;
  LPM_q_ivl_38442 <= tmp_ivl_38444 & tmp_ivl_38439;
  tmp_ivl_38447 <= fresh(114);
  LPM_q_ivl_38449 <= tmp_ivl_38451 & tmp_ivl_38447;
  new_AGEMA_signal_3569 <= tmp_ivl_38455(1);
  tmp_ivl_38453 <= tmp_ivl_38455(0);
  tmp_ivl_38455 <= LPM_d0_ivl_38459(0 + 1 downto 0);
  tmp_ivl_38461 <= y4(56);
  tmp_ivl_38462 <= new_AGEMA_signal_2374 & tmp_ivl_38461;
  LPM_q_ivl_38465 <= tmp_ivl_38467 & tmp_ivl_38462;
  tmp_ivl_38469 <= new_AGEMA_signal_3098 & SboxInst_n269;
  LPM_q_ivl_38472 <= tmp_ivl_38474 & tmp_ivl_38469;
  tmp_ivl_38477 <= fresh(115);
  LPM_q_ivl_38479 <= tmp_ivl_38481 & tmp_ivl_38477;
  new_AGEMA_signal_3570 <= tmp_ivl_38485(1);
  tmp_ivl_38483 <= tmp_ivl_38485(0);
  tmp_ivl_38485 <= LPM_d0_ivl_38489(0 + 1 downto 0);
  tmp_ivl_38491 <= y4(57);
  tmp_ivl_38492 <= new_AGEMA_signal_2371 & tmp_ivl_38491;
  LPM_q_ivl_38495 <= tmp_ivl_38497 & tmp_ivl_38492;
  tmp_ivl_38499 <= new_AGEMA_signal_3099 & SboxInst_n268;
  LPM_q_ivl_38502 <= tmp_ivl_38504 & tmp_ivl_38499;
  tmp_ivl_38507 <= fresh(116);
  LPM_q_ivl_38509 <= tmp_ivl_38511 & tmp_ivl_38507;
  new_AGEMA_signal_3571 <= tmp_ivl_38515(1);
  tmp_ivl_38513 <= tmp_ivl_38515(0);
  tmp_ivl_38515 <= LPM_d0_ivl_38519(0 + 1 downto 0);
  tmp_ivl_38521 <= y4(58);
  tmp_ivl_38522 <= new_AGEMA_signal_2368 & tmp_ivl_38521;
  LPM_q_ivl_38525 <= tmp_ivl_38527 & tmp_ivl_38522;
  tmp_ivl_38529 <= new_AGEMA_signal_3100 & SboxInst_n267;
  LPM_q_ivl_38532 <= tmp_ivl_38534 & tmp_ivl_38529;
  tmp_ivl_38537 <= fresh(117);
  LPM_q_ivl_38539 <= tmp_ivl_38541 & tmp_ivl_38537;
  new_AGEMA_signal_3572 <= tmp_ivl_38545(1);
  tmp_ivl_38543 <= tmp_ivl_38545(0);
  tmp_ivl_38545 <= LPM_d0_ivl_38549(0 + 1 downto 0);
  tmp_ivl_38551 <= y4(59);
  tmp_ivl_38552 <= new_AGEMA_signal_2365 & tmp_ivl_38551;
  LPM_q_ivl_38555 <= tmp_ivl_38557 & tmp_ivl_38552;
  tmp_ivl_38559 <= new_AGEMA_signal_3101 & SboxInst_n266;
  LPM_q_ivl_38562 <= tmp_ivl_38564 & tmp_ivl_38559;
  tmp_ivl_38567 <= fresh(118);
  LPM_q_ivl_38569 <= tmp_ivl_38571 & tmp_ivl_38567;
  new_AGEMA_signal_3573 <= tmp_ivl_38575(1);
  tmp_ivl_38573 <= tmp_ivl_38575(0);
  tmp_ivl_38575 <= LPM_d0_ivl_38579(0 + 1 downto 0);
  tmp_ivl_38581 <= y4(5);
  tmp_ivl_38582 <= new_AGEMA_signal_2362 & tmp_ivl_38581;
  LPM_q_ivl_38585 <= tmp_ivl_38587 & tmp_ivl_38582;
  tmp_ivl_38589 <= new_AGEMA_signal_3102 & SboxInst_n265;
  LPM_q_ivl_38592 <= tmp_ivl_38594 & tmp_ivl_38589;
  tmp_ivl_38597 <= fresh(119);
  LPM_q_ivl_38599 <= tmp_ivl_38601 & tmp_ivl_38597;
  new_AGEMA_signal_3574 <= tmp_ivl_38605(1);
  tmp_ivl_38603 <= tmp_ivl_38605(0);
  tmp_ivl_38605 <= LPM_d0_ivl_38609(0 + 1 downto 0);
  tmp_ivl_38611 <= y4(60);
  tmp_ivl_38612 <= new_AGEMA_signal_2359 & tmp_ivl_38611;
  LPM_q_ivl_38615 <= tmp_ivl_38617 & tmp_ivl_38612;
  tmp_ivl_38619 <= new_AGEMA_signal_3103 & SboxInst_n264;
  LPM_q_ivl_38622 <= tmp_ivl_38624 & tmp_ivl_38619;
  tmp_ivl_38627 <= fresh(120);
  LPM_q_ivl_38629 <= tmp_ivl_38631 & tmp_ivl_38627;
  new_AGEMA_signal_3575 <= tmp_ivl_38635(1);
  tmp_ivl_38633 <= tmp_ivl_38635(0);
  tmp_ivl_38635 <= LPM_d0_ivl_38639(0 + 1 downto 0);
  tmp_ivl_38641 <= y4(61);
  tmp_ivl_38642 <= new_AGEMA_signal_2356 & tmp_ivl_38641;
  LPM_q_ivl_38645 <= tmp_ivl_38647 & tmp_ivl_38642;
  tmp_ivl_38649 <= new_AGEMA_signal_3104 & SboxInst_n263;
  LPM_q_ivl_38652 <= tmp_ivl_38654 & tmp_ivl_38649;
  tmp_ivl_38657 <= fresh(121);
  LPM_q_ivl_38659 <= tmp_ivl_38661 & tmp_ivl_38657;
  new_AGEMA_signal_3576 <= tmp_ivl_38665(1);
  tmp_ivl_38663 <= tmp_ivl_38665(0);
  tmp_ivl_38665 <= LPM_d0_ivl_38669(0 + 1 downto 0);
  tmp_ivl_38671 <= y4(62);
  tmp_ivl_38672 <= new_AGEMA_signal_2353 & tmp_ivl_38671;
  LPM_q_ivl_38675 <= tmp_ivl_38677 & tmp_ivl_38672;
  tmp_ivl_38679 <= new_AGEMA_signal_3105 & SboxInst_n262;
  LPM_q_ivl_38682 <= tmp_ivl_38684 & tmp_ivl_38679;
  tmp_ivl_38687 <= fresh(122);
  LPM_q_ivl_38689 <= tmp_ivl_38691 & tmp_ivl_38687;
  new_AGEMA_signal_3577 <= tmp_ivl_38695(1);
  tmp_ivl_38693 <= tmp_ivl_38695(0);
  tmp_ivl_38695 <= LPM_d0_ivl_38699(0 + 1 downto 0);
  tmp_ivl_38701 <= y4(63);
  tmp_ivl_38702 <= new_AGEMA_signal_2350 & tmp_ivl_38701;
  LPM_q_ivl_38705 <= tmp_ivl_38707 & tmp_ivl_38702;
  tmp_ivl_38709 <= new_AGEMA_signal_3106 & SboxInst_n261;
  LPM_q_ivl_38712 <= tmp_ivl_38714 & tmp_ivl_38709;
  tmp_ivl_38717 <= fresh(123);
  LPM_q_ivl_38719 <= tmp_ivl_38721 & tmp_ivl_38717;
  new_AGEMA_signal_3578 <= tmp_ivl_38725(1);
  tmp_ivl_38723 <= tmp_ivl_38725(0);
  tmp_ivl_38725 <= LPM_d0_ivl_38729(0 + 1 downto 0);
  tmp_ivl_38731 <= y4(6);
  tmp_ivl_38732 <= new_AGEMA_signal_2347 & tmp_ivl_38731;
  LPM_q_ivl_38735 <= tmp_ivl_38737 & tmp_ivl_38732;
  tmp_ivl_38739 <= new_AGEMA_signal_3107 & SboxInst_n260;
  LPM_q_ivl_38742 <= tmp_ivl_38744 & tmp_ivl_38739;
  tmp_ivl_38747 <= fresh(124);
  LPM_q_ivl_38749 <= tmp_ivl_38751 & tmp_ivl_38747;
  new_AGEMA_signal_3579 <= tmp_ivl_38755(1);
  tmp_ivl_38753 <= tmp_ivl_38755(0);
  tmp_ivl_38755 <= LPM_d0_ivl_38759(0 + 1 downto 0);
  tmp_ivl_38761 <= y4(7);
  tmp_ivl_38762 <= new_AGEMA_signal_2344 & tmp_ivl_38761;
  LPM_q_ivl_38765 <= tmp_ivl_38767 & tmp_ivl_38762;
  tmp_ivl_38769 <= new_AGEMA_signal_3108 & SboxInst_n259;
  LPM_q_ivl_38772 <= tmp_ivl_38774 & tmp_ivl_38769;
  tmp_ivl_38777 <= fresh(125);
  LPM_q_ivl_38779 <= tmp_ivl_38781 & tmp_ivl_38777;
  new_AGEMA_signal_3580 <= tmp_ivl_38785(1);
  tmp_ivl_38783 <= tmp_ivl_38785(0);
  tmp_ivl_38785 <= LPM_d0_ivl_38789(0 + 1 downto 0);
  tmp_ivl_38791 <= y4(8);
  tmp_ivl_38792 <= new_AGEMA_signal_2341 & tmp_ivl_38791;
  LPM_q_ivl_38795 <= tmp_ivl_38797 & tmp_ivl_38792;
  tmp_ivl_38799 <= new_AGEMA_signal_3109 & SboxInst_n258;
  LPM_q_ivl_38802 <= tmp_ivl_38804 & tmp_ivl_38799;
  tmp_ivl_38807 <= fresh(126);
  LPM_q_ivl_38809 <= tmp_ivl_38811 & tmp_ivl_38807;
  new_AGEMA_signal_3581 <= tmp_ivl_38815(1);
  tmp_ivl_38813 <= tmp_ivl_38815(0);
  tmp_ivl_38815 <= LPM_d0_ivl_38819(0 + 1 downto 0);
  tmp_ivl_38821 <= y4(9);
  tmp_ivl_38822 <= new_AGEMA_signal_2338 & tmp_ivl_38821;
  LPM_q_ivl_38825 <= tmp_ivl_38827 & tmp_ivl_38822;
  tmp_ivl_38829 <= new_AGEMA_signal_3110 & SboxInst_n257;
  LPM_q_ivl_38832 <= tmp_ivl_38834 & tmp_ivl_38829;
  tmp_ivl_38837 <= fresh(127);
  LPM_q_ivl_38839 <= tmp_ivl_38841 & tmp_ivl_38837;
  new_AGEMA_signal_3582 <= tmp_ivl_38845(1);
  tmp_ivl_38843 <= tmp_ivl_38845(0);
  tmp_ivl_38845 <= LPM_d0_ivl_38849(0 + 1 downto 0);
  tmp_ivl_38851 <= y0(0);
  tmp_ivl_38852 <= new_AGEMA_signal_2655 & tmp_ivl_38851;
  LPM_q_ivl_38855 <= tmp_ivl_38857 & tmp_ivl_38852;
  tmp_ivl_38859 <= new_AGEMA_signal_2911 & SboxInst_n256;
  LPM_q_ivl_38862 <= tmp_ivl_38864 & tmp_ivl_38859;
  tmp_ivl_38867 <= fresh(128);
  LPM_q_ivl_38869 <= tmp_ivl_38871 & tmp_ivl_38867;
  new_AGEMA_signal_3111 <= tmp_ivl_38875(1);
  tmp_ivl_38873 <= tmp_ivl_38875(0);
  tmp_ivl_38875 <= LPM_d0_ivl_38879(0 + 1 downto 0);
  tmp_ivl_38881 <= y0(10);
  tmp_ivl_38882 <= new_AGEMA_signal_2653 & tmp_ivl_38881;
  LPM_q_ivl_38885 <= tmp_ivl_38887 & tmp_ivl_38882;
  tmp_ivl_38889 <= new_AGEMA_signal_2924 & SboxInst_n255;
  LPM_q_ivl_38892 <= tmp_ivl_38894 & tmp_ivl_38889;
  tmp_ivl_38897 <= fresh(129);
  LPM_q_ivl_38899 <= tmp_ivl_38901 & tmp_ivl_38897;
  new_AGEMA_signal_3112 <= tmp_ivl_38905(1);
  tmp_ivl_38903 <= tmp_ivl_38905(0);
  tmp_ivl_38905 <= LPM_d0_ivl_38909(0 + 1 downto 0);
  tmp_ivl_38911 <= y0(11);
  tmp_ivl_38912 <= new_AGEMA_signal_2651 & tmp_ivl_38911;
  LPM_q_ivl_38915 <= tmp_ivl_38917 & tmp_ivl_38912;
  tmp_ivl_38919 <= new_AGEMA_signal_2921 & SboxInst_n254;
  LPM_q_ivl_38922 <= tmp_ivl_38924 & tmp_ivl_38919;
  tmp_ivl_38927 <= fresh(130);
  LPM_q_ivl_38929 <= tmp_ivl_38931 & tmp_ivl_38927;
  new_AGEMA_signal_3113 <= tmp_ivl_38935(1);
  tmp_ivl_38933 <= tmp_ivl_38935(0);
  tmp_ivl_38935 <= LPM_d0_ivl_38939(0 + 1 downto 0);
  tmp_ivl_38941 <= y0(12);
  tmp_ivl_38942 <= new_AGEMA_signal_2649 & tmp_ivl_38941;
  LPM_q_ivl_38945 <= tmp_ivl_38947 & tmp_ivl_38942;
  tmp_ivl_38949 <= new_AGEMA_signal_2919 & SboxInst_n253;
  LPM_q_ivl_38952 <= tmp_ivl_38954 & tmp_ivl_38949;
  tmp_ivl_38957 <= fresh(131);
  LPM_q_ivl_38959 <= tmp_ivl_38961 & tmp_ivl_38957;
  new_AGEMA_signal_3114 <= tmp_ivl_38965(1);
  tmp_ivl_38963 <= tmp_ivl_38965(0);
  tmp_ivl_38965 <= LPM_d0_ivl_38969(0 + 1 downto 0);
  tmp_ivl_38971 <= y0(13);
  tmp_ivl_38972 <= new_AGEMA_signal_2647 & tmp_ivl_38971;
  LPM_q_ivl_38975 <= tmp_ivl_38977 & tmp_ivl_38972;
  tmp_ivl_38979 <= new_AGEMA_signal_2925 & SboxInst_n252;
  LPM_q_ivl_38982 <= tmp_ivl_38984 & tmp_ivl_38979;
  tmp_ivl_38987 <= fresh(132);
  LPM_q_ivl_38989 <= tmp_ivl_38991 & tmp_ivl_38987;
  new_AGEMA_signal_3115 <= tmp_ivl_38995(1);
  tmp_ivl_38993 <= tmp_ivl_38995(0);
  tmp_ivl_38995 <= LPM_d0_ivl_38999(0 + 1 downto 0);
  tmp_ivl_39001 <= y0(14);
  tmp_ivl_39002 <= new_AGEMA_signal_2645 & tmp_ivl_39001;
  LPM_q_ivl_39005 <= tmp_ivl_39007 & tmp_ivl_39002;
  tmp_ivl_39009 <= new_AGEMA_signal_2922 & SboxInst_n251;
  LPM_q_ivl_39012 <= tmp_ivl_39014 & tmp_ivl_39009;
  tmp_ivl_39017 <= fresh(133);
  LPM_q_ivl_39019 <= tmp_ivl_39021 & tmp_ivl_39017;
  new_AGEMA_signal_3116 <= tmp_ivl_39025(1);
  tmp_ivl_39023 <= tmp_ivl_39025(0);
  tmp_ivl_39025 <= LPM_d0_ivl_39029(0 + 1 downto 0);
  tmp_ivl_39031 <= y0(15);
  tmp_ivl_39032 <= new_AGEMA_signal_2643 & tmp_ivl_39031;
  LPM_q_ivl_39035 <= tmp_ivl_39037 & tmp_ivl_39032;
  tmp_ivl_39039 <= new_AGEMA_signal_2918 & SboxInst_n250;
  LPM_q_ivl_39042 <= tmp_ivl_39044 & tmp_ivl_39039;
  tmp_ivl_39047 <= fresh(134);
  LPM_q_ivl_39049 <= tmp_ivl_39051 & tmp_ivl_39047;
  new_AGEMA_signal_3117 <= tmp_ivl_39055(1);
  tmp_ivl_39053 <= tmp_ivl_39055(0);
  tmp_ivl_39055 <= LPM_d0_ivl_39059(0 + 1 downto 0);
  tmp_ivl_39061 <= y0(16);
  tmp_ivl_39062 <= new_AGEMA_signal_2641 & tmp_ivl_39061;
  LPM_q_ivl_39065 <= tmp_ivl_39067 & tmp_ivl_39062;
  tmp_ivl_39069 <= new_AGEMA_signal_2944 & SboxInst_n249;
  LPM_q_ivl_39072 <= tmp_ivl_39074 & tmp_ivl_39069;
  tmp_ivl_39077 <= fresh(135);
  LPM_q_ivl_39079 <= tmp_ivl_39081 & tmp_ivl_39077;
  new_AGEMA_signal_3118 <= tmp_ivl_39085(1);
  tmp_ivl_39083 <= tmp_ivl_39085(0);
  tmp_ivl_39085 <= LPM_d0_ivl_39089(0 + 1 downto 0);
  tmp_ivl_39091 <= y0(17);
  tmp_ivl_39092 <= new_AGEMA_signal_2639 & tmp_ivl_39091;
  LPM_q_ivl_39095 <= tmp_ivl_39097 & tmp_ivl_39092;
  tmp_ivl_39099 <= new_AGEMA_signal_2942 & SboxInst_n248;
  LPM_q_ivl_39102 <= tmp_ivl_39104 & tmp_ivl_39099;
  tmp_ivl_39107 <= fresh(136);
  LPM_q_ivl_39109 <= tmp_ivl_39111 & tmp_ivl_39107;
  new_AGEMA_signal_3119 <= tmp_ivl_39115(1);
  tmp_ivl_39113 <= tmp_ivl_39115(0);
  tmp_ivl_39115 <= LPM_d0_ivl_39119(0 + 1 downto 0);
  tmp_ivl_39121 <= y0(18);
  tmp_ivl_39122 <= new_AGEMA_signal_2637 & tmp_ivl_39121;
  LPM_q_ivl_39125 <= tmp_ivl_39127 & tmp_ivl_39122;
  tmp_ivl_39129 <= new_AGEMA_signal_2940 & SboxInst_n247;
  LPM_q_ivl_39132 <= tmp_ivl_39134 & tmp_ivl_39129;
  tmp_ivl_39137 <= fresh(137);
  LPM_q_ivl_39139 <= tmp_ivl_39141 & tmp_ivl_39137;
  new_AGEMA_signal_3120 <= tmp_ivl_39145(1);
  tmp_ivl_39143 <= tmp_ivl_39145(0);
  tmp_ivl_39145 <= LPM_d0_ivl_39149(0 + 1 downto 0);
  tmp_ivl_39151 <= y0(19);
  tmp_ivl_39152 <= new_AGEMA_signal_2635 & tmp_ivl_39151;
  LPM_q_ivl_39155 <= tmp_ivl_39157 & tmp_ivl_39152;
  tmp_ivl_39159 <= new_AGEMA_signal_2936 & SboxInst_n246;
  LPM_q_ivl_39162 <= tmp_ivl_39164 & tmp_ivl_39159;
  tmp_ivl_39167 <= fresh(138);
  LPM_q_ivl_39169 <= tmp_ivl_39171 & tmp_ivl_39167;
  new_AGEMA_signal_3121 <= tmp_ivl_39175(1);
  tmp_ivl_39173 <= tmp_ivl_39175(0);
  tmp_ivl_39175 <= LPM_d0_ivl_39179(0 + 1 downto 0);
  tmp_ivl_39181 <= y0(1);
  tmp_ivl_39182 <= new_AGEMA_signal_2633 & tmp_ivl_39181;
  LPM_q_ivl_39185 <= tmp_ivl_39187 & tmp_ivl_39182;
  tmp_ivl_39189 <= new_AGEMA_signal_2909 & SboxInst_n245;
  LPM_q_ivl_39192 <= tmp_ivl_39194 & tmp_ivl_39189;
  tmp_ivl_39197 <= fresh(139);
  LPM_q_ivl_39199 <= tmp_ivl_39201 & tmp_ivl_39197;
  new_AGEMA_signal_3122 <= tmp_ivl_39205(1);
  tmp_ivl_39203 <= tmp_ivl_39205(0);
  tmp_ivl_39205 <= LPM_d0_ivl_39209(0 + 1 downto 0);
  tmp_ivl_39211 <= y0(20);
  tmp_ivl_39212 <= new_AGEMA_signal_2631 & tmp_ivl_39211;
  LPM_q_ivl_39215 <= tmp_ivl_39217 & tmp_ivl_39212;
  tmp_ivl_39219 <= new_AGEMA_signal_2934 & SboxInst_n244;
  LPM_q_ivl_39222 <= tmp_ivl_39224 & tmp_ivl_39219;
  tmp_ivl_39227 <= fresh(140);
  LPM_q_ivl_39229 <= tmp_ivl_39231 & tmp_ivl_39227;
  new_AGEMA_signal_3123 <= tmp_ivl_39235(1);
  tmp_ivl_39233 <= tmp_ivl_39235(0);
  tmp_ivl_39235 <= LPM_d0_ivl_39239(0 + 1 downto 0);
  tmp_ivl_39241 <= y0(21);
  tmp_ivl_39242 <= new_AGEMA_signal_2629 & tmp_ivl_39241;
  LPM_q_ivl_39245 <= tmp_ivl_39247 & tmp_ivl_39242;
  tmp_ivl_39249 <= new_AGEMA_signal_2939 & SboxInst_n243;
  LPM_q_ivl_39252 <= tmp_ivl_39254 & tmp_ivl_39249;
  tmp_ivl_39257 <= fresh(141);
  LPM_q_ivl_39259 <= tmp_ivl_39261 & tmp_ivl_39257;
  new_AGEMA_signal_3124 <= tmp_ivl_39265(1);
  tmp_ivl_39263 <= tmp_ivl_39265(0);
  tmp_ivl_39265 <= LPM_d0_ivl_39269(0 + 1 downto 0);
  tmp_ivl_39271 <= y0(22);
  tmp_ivl_39272 <= new_AGEMA_signal_2627 & tmp_ivl_39271;
  LPM_q_ivl_39275 <= tmp_ivl_39277 & tmp_ivl_39272;
  tmp_ivl_39279 <= new_AGEMA_signal_2937 & SboxInst_n242;
  LPM_q_ivl_39282 <= tmp_ivl_39284 & tmp_ivl_39279;
  tmp_ivl_39287 <= fresh(142);
  LPM_q_ivl_39289 <= tmp_ivl_39291 & tmp_ivl_39287;
  new_AGEMA_signal_3125 <= tmp_ivl_39295(1);
  tmp_ivl_39293 <= tmp_ivl_39295(0);
  tmp_ivl_39295 <= LPM_d0_ivl_39299(0 + 1 downto 0);
  tmp_ivl_39301 <= y0(23);
  tmp_ivl_39302 <= new_AGEMA_signal_2625 & tmp_ivl_39301;
  LPM_q_ivl_39305 <= tmp_ivl_39307 & tmp_ivl_39302;
  tmp_ivl_39309 <= new_AGEMA_signal_2935 & SboxInst_n241;
  LPM_q_ivl_39312 <= tmp_ivl_39314 & tmp_ivl_39309;
  tmp_ivl_39317 <= fresh(143);
  LPM_q_ivl_39319 <= tmp_ivl_39321 & tmp_ivl_39317;
  new_AGEMA_signal_3126 <= tmp_ivl_39325(1);
  tmp_ivl_39323 <= tmp_ivl_39325(0);
  tmp_ivl_39325 <= LPM_d0_ivl_39329(0 + 1 downto 0);
  tmp_ivl_39331 <= y0(24);
  tmp_ivl_39332 <= new_AGEMA_signal_2623 & tmp_ivl_39331;
  LPM_q_ivl_39335 <= tmp_ivl_39337 & tmp_ivl_39332;
  tmp_ivl_39339 <= new_AGEMA_signal_2955 & SboxInst_n240;
  LPM_q_ivl_39342 <= tmp_ivl_39344 & tmp_ivl_39339;
  tmp_ivl_39347 <= fresh(144);
  LPM_q_ivl_39349 <= tmp_ivl_39351 & tmp_ivl_39347;
  new_AGEMA_signal_3127 <= tmp_ivl_39355(1);
  tmp_ivl_39353 <= tmp_ivl_39355(0);
  tmp_ivl_39355 <= LPM_d0_ivl_39359(0 + 1 downto 0);
  tmp_ivl_39361 <= y0(25);
  tmp_ivl_39362 <= new_AGEMA_signal_2621 & tmp_ivl_39361;
  LPM_q_ivl_39365 <= tmp_ivl_39367 & tmp_ivl_39362;
  tmp_ivl_39369 <= new_AGEMA_signal_2954 & SboxInst_n239;
  LPM_q_ivl_39372 <= tmp_ivl_39374 & tmp_ivl_39369;
  tmp_ivl_39377 <= fresh(145);
  LPM_q_ivl_39379 <= tmp_ivl_39381 & tmp_ivl_39377;
  new_AGEMA_signal_3128 <= tmp_ivl_39385(1);
  tmp_ivl_39383 <= tmp_ivl_39385(0);
  tmp_ivl_39385 <= LPM_d0_ivl_39389(0 + 1 downto 0);
  tmp_ivl_39391 <= y0(26);
  tmp_ivl_39392 <= new_AGEMA_signal_2619 & tmp_ivl_39391;
  LPM_q_ivl_39395 <= tmp_ivl_39397 & tmp_ivl_39392;
  tmp_ivl_39399 <= new_AGEMA_signal_2952 & SboxInst_n238;
  LPM_q_ivl_39402 <= tmp_ivl_39404 & tmp_ivl_39399;
  tmp_ivl_39407 <= fresh(146);
  LPM_q_ivl_39409 <= tmp_ivl_39411 & tmp_ivl_39407;
  new_AGEMA_signal_3129 <= tmp_ivl_39415(1);
  tmp_ivl_39413 <= tmp_ivl_39415(0);
  tmp_ivl_39415 <= LPM_d0_ivl_39419(0 + 1 downto 0);
  tmp_ivl_39421 <= y0(27);
  tmp_ivl_39422 <= new_AGEMA_signal_2617 & tmp_ivl_39421;
  LPM_q_ivl_39425 <= tmp_ivl_39427 & tmp_ivl_39422;
  tmp_ivl_39429 <= new_AGEMA_signal_2951 & SboxInst_n237;
  LPM_q_ivl_39432 <= tmp_ivl_39434 & tmp_ivl_39429;
  tmp_ivl_39437 <= fresh(147);
  LPM_q_ivl_39439 <= tmp_ivl_39441 & tmp_ivl_39437;
  new_AGEMA_signal_3130 <= tmp_ivl_39445(1);
  tmp_ivl_39443 <= tmp_ivl_39445(0);
  tmp_ivl_39445 <= LPM_d0_ivl_39449(0 + 1 downto 0);
  tmp_ivl_39451 <= y0(28);
  tmp_ivl_39452 <= new_AGEMA_signal_2615 & tmp_ivl_39451;
  LPM_q_ivl_39455 <= tmp_ivl_39457 & tmp_ivl_39452;
  tmp_ivl_39459 <= new_AGEMA_signal_2949 & SboxInst_n236;
  LPM_q_ivl_39462 <= tmp_ivl_39464 & tmp_ivl_39459;
  tmp_ivl_39467 <= fresh(148);
  LPM_q_ivl_39469 <= tmp_ivl_39471 & tmp_ivl_39467;
  new_AGEMA_signal_3131 <= tmp_ivl_39475(1);
  tmp_ivl_39473 <= tmp_ivl_39475(0);
  tmp_ivl_39475 <= LPM_d0_ivl_39479(0 + 1 downto 0);
  tmp_ivl_39481 <= y0(29);
  tmp_ivl_39482 <= new_AGEMA_signal_2613 & tmp_ivl_39481;
  LPM_q_ivl_39485 <= tmp_ivl_39487 & tmp_ivl_39482;
  tmp_ivl_39489 <= new_AGEMA_signal_2953 & SboxInst_n235;
  LPM_q_ivl_39492 <= tmp_ivl_39494 & tmp_ivl_39489;
  tmp_ivl_39497 <= fresh(149);
  LPM_q_ivl_39499 <= tmp_ivl_39501 & tmp_ivl_39497;
  new_AGEMA_signal_3132 <= tmp_ivl_39505(1);
  tmp_ivl_39503 <= tmp_ivl_39505(0);
  tmp_ivl_39505 <= LPM_d0_ivl_39509(0 + 1 downto 0);
  tmp_ivl_39511 <= y0(2);
  tmp_ivl_39512 <= new_AGEMA_signal_2611 & tmp_ivl_39511;
  LPM_q_ivl_39515 <= tmp_ivl_39517 & tmp_ivl_39512;
  tmp_ivl_39519 <= new_AGEMA_signal_2906 & SboxInst_n234;
  LPM_q_ivl_39522 <= tmp_ivl_39524 & tmp_ivl_39519;
  tmp_ivl_39527 <= fresh(150);
  LPM_q_ivl_39529 <= tmp_ivl_39531 & tmp_ivl_39527;
  new_AGEMA_signal_3133 <= tmp_ivl_39535(1);
  tmp_ivl_39533 <= tmp_ivl_39535(0);
  tmp_ivl_39535 <= LPM_d0_ivl_39539(0 + 1 downto 0);
  tmp_ivl_39541 <= y0(30);
  tmp_ivl_39542 <= new_AGEMA_signal_2609 & tmp_ivl_39541;
  LPM_q_ivl_39545 <= tmp_ivl_39547 & tmp_ivl_39542;
  tmp_ivl_39549 <= new_AGEMA_signal_2950 & SboxInst_n233;
  LPM_q_ivl_39552 <= tmp_ivl_39554 & tmp_ivl_39549;
  tmp_ivl_39557 <= fresh(151);
  LPM_q_ivl_39559 <= tmp_ivl_39561 & tmp_ivl_39557;
  new_AGEMA_signal_3134 <= tmp_ivl_39565(1);
  tmp_ivl_39563 <= tmp_ivl_39565(0);
  tmp_ivl_39565 <= LPM_d0_ivl_39569(0 + 1 downto 0);
  tmp_ivl_39571 <= y0(31);
  tmp_ivl_39572 <= new_AGEMA_signal_2607 & tmp_ivl_39571;
  LPM_q_ivl_39575 <= tmp_ivl_39577 & tmp_ivl_39572;
  tmp_ivl_39579 <= new_AGEMA_signal_2948 & SboxInst_n232;
  LPM_q_ivl_39582 <= tmp_ivl_39584 & tmp_ivl_39579;
  tmp_ivl_39587 <= fresh(152);
  LPM_q_ivl_39589 <= tmp_ivl_39591 & tmp_ivl_39587;
  new_AGEMA_signal_3135 <= tmp_ivl_39595(1);
  tmp_ivl_39593 <= tmp_ivl_39595(0);
  tmp_ivl_39595 <= LPM_d0_ivl_39599(0 + 1 downto 0);
  tmp_ivl_39601 <= y0(32);
  tmp_ivl_39602 <= new_AGEMA_signal_2605 & tmp_ivl_39601;
  LPM_q_ivl_39605 <= tmp_ivl_39607 & tmp_ivl_39602;
  tmp_ivl_39609 <= new_AGEMA_signal_2962 & SboxInst_n231;
  LPM_q_ivl_39612 <= tmp_ivl_39614 & tmp_ivl_39609;
  tmp_ivl_39617 <= fresh(153);
  LPM_q_ivl_39619 <= tmp_ivl_39621 & tmp_ivl_39617;
  new_AGEMA_signal_3136 <= tmp_ivl_39625(1);
  tmp_ivl_39623 <= tmp_ivl_39625(0);
  tmp_ivl_39625 <= LPM_d0_ivl_39629(0 + 1 downto 0);
  tmp_ivl_39631 <= y0(33);
  tmp_ivl_39632 <= new_AGEMA_signal_2603 & tmp_ivl_39631;
  LPM_q_ivl_39635 <= tmp_ivl_39637 & tmp_ivl_39632;
  tmp_ivl_39639 <= new_AGEMA_signal_2961 & SboxInst_n230;
  LPM_q_ivl_39642 <= tmp_ivl_39644 & tmp_ivl_39639;
  tmp_ivl_39647 <= fresh(154);
  LPM_q_ivl_39649 <= tmp_ivl_39651 & tmp_ivl_39647;
  new_AGEMA_signal_3137 <= tmp_ivl_39655(1);
  tmp_ivl_39653 <= tmp_ivl_39655(0);
  tmp_ivl_39655 <= LPM_d0_ivl_39659(0 + 1 downto 0);
  tmp_ivl_39661 <= y0(34);
  tmp_ivl_39662 <= new_AGEMA_signal_2601 & tmp_ivl_39661;
  LPM_q_ivl_39665 <= tmp_ivl_39667 & tmp_ivl_39662;
  tmp_ivl_39669 <= new_AGEMA_signal_2959 & SboxInst_n229;
  LPM_q_ivl_39672 <= tmp_ivl_39674 & tmp_ivl_39669;
  tmp_ivl_39677 <= fresh(155);
  LPM_q_ivl_39679 <= tmp_ivl_39681 & tmp_ivl_39677;
  new_AGEMA_signal_3138 <= tmp_ivl_39685(1);
  tmp_ivl_39683 <= tmp_ivl_39685(0);
  tmp_ivl_39685 <= LPM_d0_ivl_39689(0 + 1 downto 0);
  tmp_ivl_39691 <= y0(35);
  tmp_ivl_39692 <= new_AGEMA_signal_2599 & tmp_ivl_39691;
  LPM_q_ivl_39695 <= tmp_ivl_39697 & tmp_ivl_39692;
  tmp_ivl_39699 <= new_AGEMA_signal_2957 & SboxInst_n228;
  LPM_q_ivl_39702 <= tmp_ivl_39704 & tmp_ivl_39699;
  tmp_ivl_39707 <= fresh(156);
  LPM_q_ivl_39709 <= tmp_ivl_39711 & tmp_ivl_39707;
  new_AGEMA_signal_3139 <= tmp_ivl_39715(1);
  tmp_ivl_39713 <= tmp_ivl_39715(0);
  tmp_ivl_39715 <= LPM_d0_ivl_39719(0 + 1 downto 0);
  tmp_ivl_39721 <= y0(36);
  tmp_ivl_39722 <= new_AGEMA_signal_2597 & tmp_ivl_39721;
  LPM_q_ivl_39725 <= tmp_ivl_39727 & tmp_ivl_39722;
  tmp_ivl_39729 <= new_AGEMA_signal_2956 & SboxInst_n227;
  LPM_q_ivl_39732 <= tmp_ivl_39734 & tmp_ivl_39729;
  tmp_ivl_39737 <= fresh(157);
  LPM_q_ivl_39739 <= tmp_ivl_39741 & tmp_ivl_39737;
  new_AGEMA_signal_3140 <= tmp_ivl_39745(1);
  tmp_ivl_39743 <= tmp_ivl_39745(0);
  tmp_ivl_39745 <= LPM_d0_ivl_39749(0 + 1 downto 0);
  tmp_ivl_39751 <= y0(37);
  tmp_ivl_39752 <= new_AGEMA_signal_2595 & tmp_ivl_39751;
  LPM_q_ivl_39755 <= tmp_ivl_39757 & tmp_ivl_39752;
  tmp_ivl_39759 <= new_AGEMA_signal_2960 & SboxInst_n226;
  LPM_q_ivl_39762 <= tmp_ivl_39764 & tmp_ivl_39759;
  tmp_ivl_39767 <= fresh(158);
  LPM_q_ivl_39769 <= tmp_ivl_39771 & tmp_ivl_39767;
  new_AGEMA_signal_3141 <= tmp_ivl_39775(1);
  tmp_ivl_39773 <= tmp_ivl_39775(0);
  tmp_ivl_39775 <= LPM_d0_ivl_39779(0 + 1 downto 0);
  tmp_ivl_39781 <= y0(38);
  tmp_ivl_39782 <= new_AGEMA_signal_2593 & tmp_ivl_39781;
  LPM_q_ivl_39785 <= tmp_ivl_39787 & tmp_ivl_39782;
  tmp_ivl_39789 <= new_AGEMA_signal_2958 & SboxInst_n225;
  LPM_q_ivl_39792 <= tmp_ivl_39794 & tmp_ivl_39789;
  tmp_ivl_39797 <= fresh(159);
  LPM_q_ivl_39799 <= tmp_ivl_39801 & tmp_ivl_39797;
  new_AGEMA_signal_3142 <= tmp_ivl_39805(1);
  tmp_ivl_39803 <= tmp_ivl_39805(0);
  tmp_ivl_39805 <= LPM_d0_ivl_39809(0 + 1 downto 0);
  tmp_ivl_39811 <= y0(39);
  tmp_ivl_39812 <= new_AGEMA_signal_2591 & tmp_ivl_39811;
  LPM_q_ivl_39815 <= tmp_ivl_39817 & tmp_ivl_39812;
  tmp_ivl_39819 <= new_AGEMA_signal_2916 & SboxInst_n224;
  LPM_q_ivl_39822 <= tmp_ivl_39824 & tmp_ivl_39819;
  tmp_ivl_39827 <= fresh(160);
  LPM_q_ivl_39829 <= tmp_ivl_39831 & tmp_ivl_39827;
  new_AGEMA_signal_3143 <= tmp_ivl_39835(1);
  tmp_ivl_39833 <= tmp_ivl_39835(0);
  tmp_ivl_39835 <= LPM_d0_ivl_39839(0 + 1 downto 0);
  tmp_ivl_39841 <= y0(3);
  tmp_ivl_39842 <= new_AGEMA_signal_2589 & tmp_ivl_39841;
  LPM_q_ivl_39845 <= tmp_ivl_39847 & tmp_ivl_39842;
  tmp_ivl_39849 <= new_AGEMA_signal_2904 & SboxInst_n223;
  LPM_q_ivl_39852 <= tmp_ivl_39854 & tmp_ivl_39849;
  tmp_ivl_39857 <= fresh(161);
  LPM_q_ivl_39859 <= tmp_ivl_39861 & tmp_ivl_39857;
  new_AGEMA_signal_3144 <= tmp_ivl_39865(1);
  tmp_ivl_39863 <= tmp_ivl_39865(0);
  tmp_ivl_39865 <= LPM_d0_ivl_39869(0 + 1 downto 0);
  tmp_ivl_39871 <= y0(40);
  tmp_ivl_39872 <= new_AGEMA_signal_2587 & tmp_ivl_39871;
  LPM_q_ivl_39875 <= tmp_ivl_39877 & tmp_ivl_39872;
  tmp_ivl_39879 <= new_AGEMA_signal_2914 & SboxInst_n222;
  LPM_q_ivl_39882 <= tmp_ivl_39884 & tmp_ivl_39879;
  tmp_ivl_39887 <= fresh(162);
  LPM_q_ivl_39889 <= tmp_ivl_39891 & tmp_ivl_39887;
  new_AGEMA_signal_3145 <= tmp_ivl_39895(1);
  tmp_ivl_39893 <= tmp_ivl_39895(0);
  tmp_ivl_39895 <= LPM_d0_ivl_39899(0 + 1 downto 0);
  tmp_ivl_39901 <= y0(41);
  tmp_ivl_39902 <= new_AGEMA_signal_2585 & tmp_ivl_39901;
  LPM_q_ivl_39905 <= tmp_ivl_39907 & tmp_ivl_39902;
  tmp_ivl_39909 <= new_AGEMA_signal_2913 & SboxInst_n221;
  LPM_q_ivl_39912 <= tmp_ivl_39914 & tmp_ivl_39909;
  tmp_ivl_39917 <= fresh(163);
  LPM_q_ivl_39919 <= tmp_ivl_39921 & tmp_ivl_39917;
  new_AGEMA_signal_3146 <= tmp_ivl_39925(1);
  tmp_ivl_39923 <= tmp_ivl_39925(0);
  tmp_ivl_39925 <= LPM_d0_ivl_39929(0 + 1 downto 0);
  tmp_ivl_39931 <= y0(42);
  tmp_ivl_39932 <= new_AGEMA_signal_2583 & tmp_ivl_39931;
  LPM_q_ivl_39935 <= tmp_ivl_39937 & tmp_ivl_39932;
  tmp_ivl_39939 <= new_AGEMA_signal_2910 & SboxInst_n220;
  LPM_q_ivl_39942 <= tmp_ivl_39944 & tmp_ivl_39939;
  tmp_ivl_39947 <= fresh(164);
  LPM_q_ivl_39949 <= tmp_ivl_39951 & tmp_ivl_39947;
  new_AGEMA_signal_3147 <= tmp_ivl_39955(1);
  tmp_ivl_39953 <= tmp_ivl_39955(0);
  tmp_ivl_39955 <= LPM_d0_ivl_39959(0 + 1 downto 0);
  tmp_ivl_39961 <= y0(43);
  tmp_ivl_39962 <= new_AGEMA_signal_2581 & tmp_ivl_39961;
  LPM_q_ivl_39965 <= tmp_ivl_39967 & tmp_ivl_39962;
  tmp_ivl_39969 <= new_AGEMA_signal_2908 & SboxInst_n219;
  LPM_q_ivl_39972 <= tmp_ivl_39974 & tmp_ivl_39969;
  tmp_ivl_39977 <= fresh(165);
  LPM_q_ivl_39979 <= tmp_ivl_39981 & tmp_ivl_39977;
  new_AGEMA_signal_3148 <= tmp_ivl_39985(1);
  tmp_ivl_39983 <= tmp_ivl_39985(0);
  tmp_ivl_39985 <= LPM_d0_ivl_39989(0 + 1 downto 0);
  tmp_ivl_39991 <= y0(44);
  tmp_ivl_39992 <= new_AGEMA_signal_2579 & tmp_ivl_39991;
  LPM_q_ivl_39995 <= tmp_ivl_39997 & tmp_ivl_39992;
  tmp_ivl_39999 <= new_AGEMA_signal_2905 & SboxInst_n218;
  LPM_q_ivl_40002 <= tmp_ivl_40004 & tmp_ivl_39999;
  tmp_ivl_40007 <= fresh(166);
  LPM_q_ivl_40009 <= tmp_ivl_40011 & tmp_ivl_40007;
  new_AGEMA_signal_3149 <= tmp_ivl_40015(1);
  tmp_ivl_40013 <= tmp_ivl_40015(0);
  tmp_ivl_40015 <= LPM_d0_ivl_40019(0 + 1 downto 0);
  tmp_ivl_40021 <= y0(45);
  tmp_ivl_40022 <= new_AGEMA_signal_2577 & tmp_ivl_40021;
  LPM_q_ivl_40025 <= tmp_ivl_40027 & tmp_ivl_40022;
  tmp_ivl_40029 <= new_AGEMA_signal_2902 & SboxInst_n217;
  LPM_q_ivl_40032 <= tmp_ivl_40034 & tmp_ivl_40029;
  tmp_ivl_40037 <= fresh(167);
  LPM_q_ivl_40039 <= tmp_ivl_40041 & tmp_ivl_40037;
  new_AGEMA_signal_3150 <= tmp_ivl_40045(1);
  tmp_ivl_40043 <= tmp_ivl_40045(0);
  tmp_ivl_40045 <= LPM_d0_ivl_40049(0 + 1 downto 0);
  tmp_ivl_40051 <= y0(46);
  tmp_ivl_40052 <= new_AGEMA_signal_2575 & tmp_ivl_40051;
  LPM_q_ivl_40055 <= tmp_ivl_40057 & tmp_ivl_40052;
  tmp_ivl_40059 <= new_AGEMA_signal_2897 & SboxInst_n216;
  LPM_q_ivl_40062 <= tmp_ivl_40064 & tmp_ivl_40059;
  tmp_ivl_40067 <= fresh(168);
  LPM_q_ivl_40069 <= tmp_ivl_40071 & tmp_ivl_40067;
  new_AGEMA_signal_3151 <= tmp_ivl_40075(1);
  tmp_ivl_40073 <= tmp_ivl_40075(0);
  tmp_ivl_40075 <= LPM_d0_ivl_40079(0 + 1 downto 0);
  tmp_ivl_40081 <= y0(47);
  tmp_ivl_40082 <= new_AGEMA_signal_2573 & tmp_ivl_40081;
  LPM_q_ivl_40085 <= tmp_ivl_40087 & tmp_ivl_40082;
  tmp_ivl_40089 <= new_AGEMA_signal_2933 & SboxInst_n215;
  LPM_q_ivl_40092 <= tmp_ivl_40094 & tmp_ivl_40089;
  tmp_ivl_40097 <= fresh(169);
  LPM_q_ivl_40099 <= tmp_ivl_40101 & tmp_ivl_40097;
  new_AGEMA_signal_3152 <= tmp_ivl_40105(1);
  tmp_ivl_40103 <= tmp_ivl_40105(0);
  tmp_ivl_40105 <= LPM_d0_ivl_40109(0 + 1 downto 0);
  tmp_ivl_40111 <= y0(48);
  tmp_ivl_40112 <= new_AGEMA_signal_2571 & tmp_ivl_40111;
  LPM_q_ivl_40115 <= tmp_ivl_40117 & tmp_ivl_40112;
  tmp_ivl_40119 <= new_AGEMA_signal_2932 & SboxInst_n214;
  LPM_q_ivl_40122 <= tmp_ivl_40124 & tmp_ivl_40119;
  tmp_ivl_40127 <= fresh(170);
  LPM_q_ivl_40129 <= tmp_ivl_40131 & tmp_ivl_40127;
  new_AGEMA_signal_3153 <= tmp_ivl_40135(1);
  tmp_ivl_40133 <= tmp_ivl_40135(0);
  tmp_ivl_40135 <= LPM_d0_ivl_40139(0 + 1 downto 0);
  tmp_ivl_40141 <= y0(49);
  tmp_ivl_40142 <= new_AGEMA_signal_2569 & tmp_ivl_40141;
  LPM_q_ivl_40145 <= tmp_ivl_40147 & tmp_ivl_40142;
  tmp_ivl_40149 <= new_AGEMA_signal_2931 & SboxInst_n213;
  LPM_q_ivl_40152 <= tmp_ivl_40154 & tmp_ivl_40149;
  tmp_ivl_40157 <= fresh(171);
  LPM_q_ivl_40159 <= tmp_ivl_40161 & tmp_ivl_40157;
  new_AGEMA_signal_3154 <= tmp_ivl_40165(1);
  tmp_ivl_40163 <= tmp_ivl_40165(0);
  tmp_ivl_40165 <= LPM_d0_ivl_40169(0 + 1 downto 0);
  tmp_ivl_40171 <= y0(4);
  tmp_ivl_40172 <= new_AGEMA_signal_2567 & tmp_ivl_40171;
  LPM_q_ivl_40175 <= tmp_ivl_40177 & tmp_ivl_40172;
  tmp_ivl_40179 <= new_AGEMA_signal_2900 & SboxInst_n212;
  LPM_q_ivl_40182 <= tmp_ivl_40184 & tmp_ivl_40179;
  tmp_ivl_40187 <= fresh(172);
  LPM_q_ivl_40189 <= tmp_ivl_40191 & tmp_ivl_40187;
  new_AGEMA_signal_3155 <= tmp_ivl_40195(1);
  tmp_ivl_40193 <= tmp_ivl_40195(0);
  tmp_ivl_40195 <= LPM_d0_ivl_40199(0 + 1 downto 0);
  tmp_ivl_40201 <= y0(50);
  tmp_ivl_40202 <= new_AGEMA_signal_2565 & tmp_ivl_40201;
  LPM_q_ivl_40205 <= tmp_ivl_40207 & tmp_ivl_40202;
  tmp_ivl_40209 <= new_AGEMA_signal_2930 & SboxInst_n211;
  LPM_q_ivl_40212 <= tmp_ivl_40214 & tmp_ivl_40209;
  tmp_ivl_40217 <= fresh(173);
  LPM_q_ivl_40219 <= tmp_ivl_40221 & tmp_ivl_40217;
  new_AGEMA_signal_3156 <= tmp_ivl_40225(1);
  tmp_ivl_40223 <= tmp_ivl_40225(0);
  tmp_ivl_40225 <= LPM_d0_ivl_40229(0 + 1 downto 0);
  tmp_ivl_40231 <= y0(51);
  tmp_ivl_40232 <= new_AGEMA_signal_2563 & tmp_ivl_40231;
  LPM_q_ivl_40235 <= tmp_ivl_40237 & tmp_ivl_40232;
  tmp_ivl_40239 <= new_AGEMA_signal_2928 & SboxInst_n210;
  LPM_q_ivl_40242 <= tmp_ivl_40244 & tmp_ivl_40239;
  tmp_ivl_40247 <= fresh(174);
  LPM_q_ivl_40249 <= tmp_ivl_40251 & tmp_ivl_40247;
  new_AGEMA_signal_3157 <= tmp_ivl_40255(1);
  tmp_ivl_40253 <= tmp_ivl_40255(0);
  tmp_ivl_40255 <= LPM_d0_ivl_40259(0 + 1 downto 0);
  tmp_ivl_40261 <= y0(52);
  tmp_ivl_40262 <= new_AGEMA_signal_2561 & tmp_ivl_40261;
  LPM_q_ivl_40265 <= tmp_ivl_40267 & tmp_ivl_40262;
  tmp_ivl_40269 <= new_AGEMA_signal_2926 & SboxInst_n209;
  LPM_q_ivl_40272 <= tmp_ivl_40274 & tmp_ivl_40269;
  tmp_ivl_40277 <= fresh(175);
  LPM_q_ivl_40279 <= tmp_ivl_40281 & tmp_ivl_40277;
  new_AGEMA_signal_3158 <= tmp_ivl_40285(1);
  tmp_ivl_40283 <= tmp_ivl_40285(0);
  tmp_ivl_40285 <= LPM_d0_ivl_40289(0 + 1 downto 0);
  tmp_ivl_40291 <= y0(53);
  tmp_ivl_40292 <= new_AGEMA_signal_2559 & tmp_ivl_40291;
  LPM_q_ivl_40295 <= tmp_ivl_40297 & tmp_ivl_40292;
  tmp_ivl_40299 <= new_AGEMA_signal_2923 & SboxInst_n208;
  LPM_q_ivl_40302 <= tmp_ivl_40304 & tmp_ivl_40299;
  tmp_ivl_40307 <= fresh(176);
  LPM_q_ivl_40309 <= tmp_ivl_40311 & tmp_ivl_40307;
  new_AGEMA_signal_3159 <= tmp_ivl_40315(1);
  tmp_ivl_40313 <= tmp_ivl_40315(0);
  tmp_ivl_40315 <= LPM_d0_ivl_40319(0 + 1 downto 0);
  tmp_ivl_40321 <= y0(54);
  tmp_ivl_40322 <= new_AGEMA_signal_2557 & tmp_ivl_40321;
  LPM_q_ivl_40325 <= tmp_ivl_40327 & tmp_ivl_40322;
  tmp_ivl_40329 <= new_AGEMA_signal_2920 & SboxInst_n207;
  LPM_q_ivl_40332 <= tmp_ivl_40334 & tmp_ivl_40329;
  tmp_ivl_40337 <= fresh(177);
  LPM_q_ivl_40339 <= tmp_ivl_40341 & tmp_ivl_40337;
  new_AGEMA_signal_3160 <= tmp_ivl_40345(1);
  tmp_ivl_40343 <= tmp_ivl_40345(0);
  tmp_ivl_40345 <= LPM_d0_ivl_40349(0 + 1 downto 0);
  tmp_ivl_40351 <= y0(55);
  tmp_ivl_40352 <= new_AGEMA_signal_2555 & tmp_ivl_40351;
  LPM_q_ivl_40355 <= tmp_ivl_40357 & tmp_ivl_40352;
  tmp_ivl_40359 <= new_AGEMA_signal_2947 & SboxInst_n206;
  LPM_q_ivl_40362 <= tmp_ivl_40364 & tmp_ivl_40359;
  tmp_ivl_40367 <= fresh(178);
  LPM_q_ivl_40369 <= tmp_ivl_40371 & tmp_ivl_40367;
  new_AGEMA_signal_3161 <= tmp_ivl_40375(1);
  tmp_ivl_40373 <= tmp_ivl_40375(0);
  tmp_ivl_40375 <= LPM_d0_ivl_40379(0 + 1 downto 0);
  tmp_ivl_40381 <= y0(56);
  tmp_ivl_40382 <= new_AGEMA_signal_2553 & tmp_ivl_40381;
  LPM_q_ivl_40385 <= tmp_ivl_40387 & tmp_ivl_40382;
  tmp_ivl_40389 <= new_AGEMA_signal_2946 & SboxInst_n205;
  LPM_q_ivl_40392 <= tmp_ivl_40394 & tmp_ivl_40389;
  tmp_ivl_40397 <= fresh(179);
  LPM_q_ivl_40399 <= tmp_ivl_40401 & tmp_ivl_40397;
  new_AGEMA_signal_3162 <= tmp_ivl_40405(1);
  tmp_ivl_40403 <= tmp_ivl_40405(0);
  tmp_ivl_40405 <= LPM_d0_ivl_40409(0 + 1 downto 0);
  tmp_ivl_40411 <= y0(57);
  tmp_ivl_40412 <= new_AGEMA_signal_2551 & tmp_ivl_40411;
  LPM_q_ivl_40415 <= tmp_ivl_40417 & tmp_ivl_40412;
  tmp_ivl_40419 <= new_AGEMA_signal_2945 & SboxInst_n204;
  LPM_q_ivl_40422 <= tmp_ivl_40424 & tmp_ivl_40419;
  tmp_ivl_40427 <= fresh(180);
  LPM_q_ivl_40429 <= tmp_ivl_40431 & tmp_ivl_40427;
  new_AGEMA_signal_3163 <= tmp_ivl_40435(1);
  tmp_ivl_40433 <= tmp_ivl_40435(0);
  tmp_ivl_40435 <= LPM_d0_ivl_40439(0 + 1 downto 0);
  tmp_ivl_40441 <= y0(58);
  tmp_ivl_40442 <= new_AGEMA_signal_2549 & tmp_ivl_40441;
  LPM_q_ivl_40445 <= tmp_ivl_40447 & tmp_ivl_40442;
  tmp_ivl_40449 <= new_AGEMA_signal_2943 & SboxInst_n203;
  LPM_q_ivl_40452 <= tmp_ivl_40454 & tmp_ivl_40449;
  tmp_ivl_40457 <= fresh(181);
  LPM_q_ivl_40459 <= tmp_ivl_40461 & tmp_ivl_40457;
  new_AGEMA_signal_3164 <= tmp_ivl_40465(1);
  tmp_ivl_40463 <= tmp_ivl_40465(0);
  tmp_ivl_40465 <= LPM_d0_ivl_40469(0 + 1 downto 0);
  tmp_ivl_40471 <= y0(59);
  tmp_ivl_40472 <= new_AGEMA_signal_2547 & tmp_ivl_40471;
  LPM_q_ivl_40475 <= tmp_ivl_40477 & tmp_ivl_40472;
  tmp_ivl_40479 <= new_AGEMA_signal_2941 & SboxInst_n202;
  LPM_q_ivl_40482 <= tmp_ivl_40484 & tmp_ivl_40479;
  tmp_ivl_40487 <= fresh(182);
  LPM_q_ivl_40489 <= tmp_ivl_40491 & tmp_ivl_40487;
  new_AGEMA_signal_3165 <= tmp_ivl_40495(1);
  tmp_ivl_40493 <= tmp_ivl_40495(0);
  tmp_ivl_40495 <= LPM_d0_ivl_40499(0 + 1 downto 0);
  tmp_ivl_40501 <= y0(5);
  tmp_ivl_40502 <= new_AGEMA_signal_2545 & tmp_ivl_40501;
  LPM_q_ivl_40505 <= tmp_ivl_40507 & tmp_ivl_40502;
  tmp_ivl_40509 <= new_AGEMA_signal_2907 & SboxInst_n201;
  LPM_q_ivl_40512 <= tmp_ivl_40514 & tmp_ivl_40509;
  tmp_ivl_40517 <= fresh(183);
  LPM_q_ivl_40519 <= tmp_ivl_40521 & tmp_ivl_40517;
  new_AGEMA_signal_3166 <= tmp_ivl_40525(1);
  tmp_ivl_40523 <= tmp_ivl_40525(0);
  tmp_ivl_40525 <= LPM_d0_ivl_40529(0 + 1 downto 0);
  tmp_ivl_40531 <= y0(60);
  tmp_ivl_40532 <= new_AGEMA_signal_2543 & tmp_ivl_40531;
  LPM_q_ivl_40535 <= tmp_ivl_40537 & tmp_ivl_40532;
  tmp_ivl_40539 <= new_AGEMA_signal_2938 & SboxInst_n200;
  LPM_q_ivl_40542 <= tmp_ivl_40544 & tmp_ivl_40539;
  tmp_ivl_40547 <= fresh(184);
  LPM_q_ivl_40549 <= tmp_ivl_40551 & tmp_ivl_40547;
  new_AGEMA_signal_3167 <= tmp_ivl_40555(1);
  tmp_ivl_40553 <= tmp_ivl_40555(0);
  tmp_ivl_40555 <= LPM_d0_ivl_40559(0 + 1 downto 0);
  tmp_ivl_40561 <= y0(61);
  tmp_ivl_40562 <= new_AGEMA_signal_2541 & tmp_ivl_40561;
  LPM_q_ivl_40565 <= tmp_ivl_40567 & tmp_ivl_40562;
  tmp_ivl_40569 <= new_AGEMA_signal_2917 & SboxInst_n199;
  LPM_q_ivl_40572 <= tmp_ivl_40574 & tmp_ivl_40569;
  tmp_ivl_40577 <= fresh(185);
  LPM_q_ivl_40579 <= tmp_ivl_40581 & tmp_ivl_40577;
  new_AGEMA_signal_3168 <= tmp_ivl_40585(1);
  tmp_ivl_40583 <= tmp_ivl_40585(0);
  tmp_ivl_40585 <= LPM_d0_ivl_40589(0 + 1 downto 0);
  tmp_ivl_40591 <= y0(62);
  tmp_ivl_40592 <= new_AGEMA_signal_2539 & tmp_ivl_40591;
  LPM_q_ivl_40595 <= tmp_ivl_40597 & tmp_ivl_40592;
  tmp_ivl_40599 <= new_AGEMA_signal_2915 & SboxInst_n198;
  LPM_q_ivl_40602 <= tmp_ivl_40604 & tmp_ivl_40599;
  tmp_ivl_40607 <= fresh(186);
  LPM_q_ivl_40609 <= tmp_ivl_40611 & tmp_ivl_40607;
  new_AGEMA_signal_3169 <= tmp_ivl_40615(1);
  tmp_ivl_40613 <= tmp_ivl_40615(0);
  tmp_ivl_40615 <= LPM_d0_ivl_40619(0 + 1 downto 0);
  tmp_ivl_40621 <= y0(63);
  tmp_ivl_40622 <= new_AGEMA_signal_2537 & tmp_ivl_40621;
  LPM_q_ivl_40625 <= tmp_ivl_40627 & tmp_ivl_40622;
  tmp_ivl_40629 <= new_AGEMA_signal_2912 & SboxInst_n197;
  LPM_q_ivl_40632 <= tmp_ivl_40634 & tmp_ivl_40629;
  tmp_ivl_40637 <= fresh(187);
  LPM_q_ivl_40639 <= tmp_ivl_40641 & tmp_ivl_40637;
  new_AGEMA_signal_3170 <= tmp_ivl_40645(1);
  tmp_ivl_40643 <= tmp_ivl_40645(0);
  tmp_ivl_40645 <= LPM_d0_ivl_40649(0 + 1 downto 0);
  tmp_ivl_40651 <= y0(6);
  tmp_ivl_40652 <= new_AGEMA_signal_2535 & tmp_ivl_40651;
  LPM_q_ivl_40655 <= tmp_ivl_40657 & tmp_ivl_40652;
  tmp_ivl_40659 <= new_AGEMA_signal_2901 & SboxInst_n196;
  LPM_q_ivl_40662 <= tmp_ivl_40664 & tmp_ivl_40659;
  tmp_ivl_40667 <= fresh(188);
  LPM_q_ivl_40669 <= tmp_ivl_40671 & tmp_ivl_40667;
  new_AGEMA_signal_3171 <= tmp_ivl_40675(1);
  tmp_ivl_40673 <= tmp_ivl_40675(0);
  tmp_ivl_40675 <= LPM_d0_ivl_40679(0 + 1 downto 0);
  tmp_ivl_40681 <= y0(7);
  tmp_ivl_40682 <= new_AGEMA_signal_2533 & tmp_ivl_40681;
  LPM_q_ivl_40685 <= tmp_ivl_40687 & tmp_ivl_40682;
  tmp_ivl_40689 <= new_AGEMA_signal_2899 & SboxInst_n195;
  LPM_q_ivl_40692 <= tmp_ivl_40694 & tmp_ivl_40689;
  tmp_ivl_40697 <= fresh(189);
  LPM_q_ivl_40699 <= tmp_ivl_40701 & tmp_ivl_40697;
  new_AGEMA_signal_3172 <= tmp_ivl_40705(1);
  tmp_ivl_40703 <= tmp_ivl_40705(0);
  tmp_ivl_40705 <= LPM_d0_ivl_40709(0 + 1 downto 0);
  tmp_ivl_40711 <= y0(8);
  tmp_ivl_40712 <= new_AGEMA_signal_2531 & tmp_ivl_40711;
  LPM_q_ivl_40715 <= tmp_ivl_40717 & tmp_ivl_40712;
  tmp_ivl_40719 <= new_AGEMA_signal_2929 & SboxInst_n194;
  LPM_q_ivl_40722 <= tmp_ivl_40724 & tmp_ivl_40719;
  tmp_ivl_40727 <= fresh(190);
  LPM_q_ivl_40729 <= tmp_ivl_40731 & tmp_ivl_40727;
  new_AGEMA_signal_3173 <= tmp_ivl_40735(1);
  tmp_ivl_40733 <= tmp_ivl_40735(0);
  tmp_ivl_40735 <= LPM_d0_ivl_40739(0 + 1 downto 0);
  tmp_ivl_40741 <= y0(9);
  tmp_ivl_40742 <= new_AGEMA_signal_2529 & tmp_ivl_40741;
  LPM_q_ivl_40745 <= tmp_ivl_40747 & tmp_ivl_40742;
  tmp_ivl_40749 <= new_AGEMA_signal_2927 & SboxInst_n193;
  LPM_q_ivl_40752 <= tmp_ivl_40754 & tmp_ivl_40749;
  tmp_ivl_40757 <= fresh(191);
  LPM_q_ivl_40759 <= tmp_ivl_40761 & tmp_ivl_40757;
  new_AGEMA_signal_3174 <= tmp_ivl_40765(1);
  tmp_ivl_40763 <= tmp_ivl_40765(0);
  tmp_ivl_40765 <= LPM_d0_ivl_40769(0 + 1 downto 0);
  tmp_ivl_40770 <= new_AGEMA_signal_2859 & SboxInst_n345;
  LPM_q_ivl_40773 <= tmp_ivl_40775 & tmp_ivl_40770;
  tmp_ivl_40778 <= y4(45);
  tmp_ivl_40779 <= new_AGEMA_signal_2410 & tmp_ivl_40778;
  LPM_q_ivl_40782 <= tmp_ivl_40784 & tmp_ivl_40779;
  tmp_ivl_40787 <= fresh(192);
  LPM_q_ivl_40789 <= tmp_ivl_40791 & tmp_ivl_40787;
  new_AGEMA_signal_3175 <= tmp_ivl_40795(1);
  tmp_ivl_40793 <= tmp_ivl_40795(0);
  tmp_ivl_40795 <= LPM_d0_ivl_40799(0 + 1 downto 0);
  tmp_ivl_40800 <= new_AGEMA_signal_2860 & SboxInst_n352;
  LPM_q_ivl_40803 <= tmp_ivl_40805 & tmp_ivl_40800;
  tmp_ivl_40808 <= y4(39);
  tmp_ivl_40809 <= new_AGEMA_signal_2431 & tmp_ivl_40808;
  LPM_q_ivl_40812 <= tmp_ivl_40814 & tmp_ivl_40809;
  tmp_ivl_40817 <= fresh(193);
  LPM_q_ivl_40819 <= tmp_ivl_40821 & tmp_ivl_40817;
  new_AGEMA_signal_3176 <= tmp_ivl_40825(1);
  tmp_ivl_40823 <= tmp_ivl_40825(0);
  tmp_ivl_40825 <= LPM_d0_ivl_40829(0 + 1 downto 0);
  tmp_ivl_40830 <= new_AGEMA_signal_2861 & SboxInst_n350;
  LPM_q_ivl_40833 <= tmp_ivl_40835 & tmp_ivl_40830;
  tmp_ivl_40838 <= y4(40);
  tmp_ivl_40839 <= new_AGEMA_signal_2425 & tmp_ivl_40838;
  LPM_q_ivl_40842 <= tmp_ivl_40844 & tmp_ivl_40839;
  tmp_ivl_40847 <= fresh(194);
  LPM_q_ivl_40849 <= tmp_ivl_40851 & tmp_ivl_40847;
  new_AGEMA_signal_3177 <= tmp_ivl_40855(1);
  tmp_ivl_40853 <= tmp_ivl_40855(0);
  tmp_ivl_40855 <= LPM_d0_ivl_40859(0 + 1 downto 0);
  tmp_ivl_40860 <= new_AGEMA_signal_2862 & SboxInst_n346;
  LPM_q_ivl_40863 <= tmp_ivl_40865 & tmp_ivl_40860;
  tmp_ivl_40868 <= y4(44);
  tmp_ivl_40869 <= new_AGEMA_signal_2413 & tmp_ivl_40868;
  LPM_q_ivl_40872 <= tmp_ivl_40874 & tmp_ivl_40869;
  tmp_ivl_40877 <= fresh(195);
  LPM_q_ivl_40879 <= tmp_ivl_40881 & tmp_ivl_40877;
  new_AGEMA_signal_3178 <= tmp_ivl_40885(1);
  tmp_ivl_40883 <= tmp_ivl_40885(0);
  tmp_ivl_40885 <= LPM_d0_ivl_40889(0 + 1 downto 0);
  tmp_ivl_40890 <= new_AGEMA_signal_2863 & SboxInst_n353;
  LPM_q_ivl_40893 <= tmp_ivl_40895 & tmp_ivl_40890;
  tmp_ivl_40898 <= y4(38);
  tmp_ivl_40899 <= new_AGEMA_signal_2434 & tmp_ivl_40898;
  LPM_q_ivl_40902 <= tmp_ivl_40904 & tmp_ivl_40899;
  tmp_ivl_40907 <= fresh(196);
  LPM_q_ivl_40909 <= tmp_ivl_40911 & tmp_ivl_40907;
  new_AGEMA_signal_3179 <= tmp_ivl_40915(1);
  tmp_ivl_40913 <= tmp_ivl_40915(0);
  tmp_ivl_40915 <= LPM_d0_ivl_40919(0 + 1 downto 0);
  tmp_ivl_40920 <= new_AGEMA_signal_2864 & SboxInst_n347;
  LPM_q_ivl_40923 <= tmp_ivl_40925 & tmp_ivl_40920;
  tmp_ivl_40928 <= y4(43);
  tmp_ivl_40929 <= new_AGEMA_signal_2416 & tmp_ivl_40928;
  LPM_q_ivl_40932 <= tmp_ivl_40934 & tmp_ivl_40929;
  tmp_ivl_40937 <= fresh(197);
  LPM_q_ivl_40939 <= tmp_ivl_40941 & tmp_ivl_40937;
  new_AGEMA_signal_3180 <= tmp_ivl_40945(1);
  tmp_ivl_40943 <= tmp_ivl_40945(0);
  tmp_ivl_40945 <= LPM_d0_ivl_40949(0 + 1 downto 0);
  tmp_ivl_40950 <= new_AGEMA_signal_2865 & SboxInst_n354;
  LPM_q_ivl_40953 <= tmp_ivl_40955 & tmp_ivl_40950;
  tmp_ivl_40958 <= y4(37);
  tmp_ivl_40959 <= new_AGEMA_signal_2437 & tmp_ivl_40958;
  LPM_q_ivl_40962 <= tmp_ivl_40964 & tmp_ivl_40959;
  tmp_ivl_40967 <= fresh(198);
  LPM_q_ivl_40969 <= tmp_ivl_40971 & tmp_ivl_40967;
  new_AGEMA_signal_3181 <= tmp_ivl_40975(1);
  tmp_ivl_40973 <= tmp_ivl_40975(0);
  tmp_ivl_40975 <= LPM_d0_ivl_40979(0 + 1 downto 0);
  tmp_ivl_40980 <= new_AGEMA_signal_2866 & SboxInst_n348;
  LPM_q_ivl_40983 <= tmp_ivl_40985 & tmp_ivl_40980;
  tmp_ivl_40988 <= y4(42);
  tmp_ivl_40989 <= new_AGEMA_signal_2419 & tmp_ivl_40988;
  LPM_q_ivl_40992 <= tmp_ivl_40994 & tmp_ivl_40989;
  tmp_ivl_40997 <= fresh(199);
  LPM_q_ivl_40999 <= tmp_ivl_41001 & tmp_ivl_40997;
  new_AGEMA_signal_3182 <= tmp_ivl_41005(1);
  tmp_ivl_41003 <= tmp_ivl_41005(0);
  tmp_ivl_41005 <= LPM_d0_ivl_41009(0 + 1 downto 0);
  tmp_ivl_41010 <= new_AGEMA_signal_2867 & SboxInst_n355;
  LPM_q_ivl_41013 <= tmp_ivl_41015 & tmp_ivl_41010;
  tmp_ivl_41018 <= y4(36);
  tmp_ivl_41019 <= new_AGEMA_signal_2440 & tmp_ivl_41018;
  LPM_q_ivl_41022 <= tmp_ivl_41024 & tmp_ivl_41019;
  tmp_ivl_41027 <= fresh(200);
  LPM_q_ivl_41029 <= tmp_ivl_41031 & tmp_ivl_41027;
  new_AGEMA_signal_3183 <= tmp_ivl_41035(1);
  tmp_ivl_41033 <= tmp_ivl_41035(0);
  tmp_ivl_41035 <= LPM_d0_ivl_41039(0 + 1 downto 0);
  tmp_ivl_41040 <= new_AGEMA_signal_2868 & SboxInst_n349;
  LPM_q_ivl_41043 <= tmp_ivl_41045 & tmp_ivl_41040;
  tmp_ivl_41048 <= y4(41);
  tmp_ivl_41049 <= new_AGEMA_signal_2422 & tmp_ivl_41048;
  LPM_q_ivl_41052 <= tmp_ivl_41054 & tmp_ivl_41049;
  tmp_ivl_41057 <= fresh(201);
  LPM_q_ivl_41059 <= tmp_ivl_41061 & tmp_ivl_41057;
  new_AGEMA_signal_3184 <= tmp_ivl_41065(1);
  tmp_ivl_41063 <= tmp_ivl_41065(0);
  tmp_ivl_41065 <= LPM_d0_ivl_41069(0 + 1 downto 0);
  tmp_ivl_41070 <= new_AGEMA_signal_2869 & SboxInst_n356;
  LPM_q_ivl_41073 <= tmp_ivl_41075 & tmp_ivl_41070;
  tmp_ivl_41078 <= y4(35);
  tmp_ivl_41079 <= new_AGEMA_signal_2443 & tmp_ivl_41078;
  LPM_q_ivl_41082 <= tmp_ivl_41084 & tmp_ivl_41079;
  tmp_ivl_41087 <= fresh(202);
  LPM_q_ivl_41089 <= tmp_ivl_41091 & tmp_ivl_41087;
  new_AGEMA_signal_3185 <= tmp_ivl_41095(1);
  tmp_ivl_41093 <= tmp_ivl_41095(0);
  tmp_ivl_41095 <= LPM_d0_ivl_41099(0 + 1 downto 0);
  tmp_ivl_41100 <= new_AGEMA_signal_2870 & SboxInst_n357;
  LPM_q_ivl_41103 <= tmp_ivl_41105 & tmp_ivl_41100;
  tmp_ivl_41108 <= y4(34);
  tmp_ivl_41109 <= new_AGEMA_signal_2446 & tmp_ivl_41108;
  LPM_q_ivl_41112 <= tmp_ivl_41114 & tmp_ivl_41109;
  tmp_ivl_41117 <= fresh(203);
  LPM_q_ivl_41119 <= tmp_ivl_41121 & tmp_ivl_41117;
  new_AGEMA_signal_3186 <= tmp_ivl_41125(1);
  tmp_ivl_41123 <= tmp_ivl_41125(0);
  tmp_ivl_41125 <= LPM_d0_ivl_41129(0 + 1 downto 0);
  tmp_ivl_41130 <= new_AGEMA_signal_2871 & SboxInst_n358;
  LPM_q_ivl_41133 <= tmp_ivl_41135 & tmp_ivl_41130;
  tmp_ivl_41138 <= y4(33);
  tmp_ivl_41139 <= new_AGEMA_signal_2449 & tmp_ivl_41138;
  LPM_q_ivl_41142 <= tmp_ivl_41144 & tmp_ivl_41139;
  tmp_ivl_41147 <= fresh(204);
  LPM_q_ivl_41149 <= tmp_ivl_41151 & tmp_ivl_41147;
  new_AGEMA_signal_3187 <= tmp_ivl_41155(1);
  tmp_ivl_41153 <= tmp_ivl_41155(0);
  tmp_ivl_41155 <= LPM_d0_ivl_41159(0 + 1 downto 0);
  tmp_ivl_41160 <= new_AGEMA_signal_2872 & SboxInst_n359;
  LPM_q_ivl_41163 <= tmp_ivl_41165 & tmp_ivl_41160;
  tmp_ivl_41168 <= y4(32);
  tmp_ivl_41169 <= new_AGEMA_signal_2452 & tmp_ivl_41168;
  LPM_q_ivl_41172 <= tmp_ivl_41174 & tmp_ivl_41169;
  tmp_ivl_41177 <= fresh(205);
  LPM_q_ivl_41179 <= tmp_ivl_41181 & tmp_ivl_41177;
  new_AGEMA_signal_3188 <= tmp_ivl_41185(1);
  tmp_ivl_41183 <= tmp_ivl_41185(0);
  tmp_ivl_41185 <= LPM_d0_ivl_41189(0 + 1 downto 0);
  tmp_ivl_41190 <= new_AGEMA_signal_2873 & SboxInst_n342;
  LPM_q_ivl_41193 <= tmp_ivl_41195 & tmp_ivl_41190;
  tmp_ivl_41198 <= y4(48);
  tmp_ivl_41199 <= new_AGEMA_signal_2401 & tmp_ivl_41198;
  LPM_q_ivl_41202 <= tmp_ivl_41204 & tmp_ivl_41199;
  tmp_ivl_41207 <= fresh(206);
  LPM_q_ivl_41209 <= tmp_ivl_41211 & tmp_ivl_41207;
  new_AGEMA_signal_3189 <= tmp_ivl_41215(1);
  tmp_ivl_41213 <= tmp_ivl_41215(0);
  tmp_ivl_41215 <= LPM_d0_ivl_41219(0 + 1 downto 0);
  tmp_ivl_41220 <= new_AGEMA_signal_2874 & SboxInst_n336;
  LPM_q_ivl_41223 <= tmp_ivl_41225 & tmp_ivl_41220;
  tmp_ivl_41228 <= y4(53);
  tmp_ivl_41229 <= new_AGEMA_signal_2383 & tmp_ivl_41228;
  LPM_q_ivl_41232 <= tmp_ivl_41234 & tmp_ivl_41229;
  tmp_ivl_41237 <= fresh(207);
  LPM_q_ivl_41239 <= tmp_ivl_41241 & tmp_ivl_41237;
  new_AGEMA_signal_3190 <= tmp_ivl_41245(1);
  tmp_ivl_41243 <= tmp_ivl_41245(0);
  tmp_ivl_41245 <= LPM_d0_ivl_41249(0 + 1 downto 0);
  tmp_ivl_41250 <= new_AGEMA_signal_2875 & SboxInst_n343;
  LPM_q_ivl_41253 <= tmp_ivl_41255 & tmp_ivl_41250;
  tmp_ivl_41258 <= y4(47);
  tmp_ivl_41259 <= new_AGEMA_signal_2404 & tmp_ivl_41258;
  LPM_q_ivl_41262 <= tmp_ivl_41264 & tmp_ivl_41259;
  tmp_ivl_41267 <= fresh(208);
  LPM_q_ivl_41269 <= tmp_ivl_41271 & tmp_ivl_41267;
  new_AGEMA_signal_3191 <= tmp_ivl_41275(1);
  tmp_ivl_41273 <= tmp_ivl_41275(0);
  tmp_ivl_41275 <= LPM_d0_ivl_41279(0 + 1 downto 0);
  tmp_ivl_41280 <= new_AGEMA_signal_2876 & SboxInst_n337;
  LPM_q_ivl_41283 <= tmp_ivl_41285 & tmp_ivl_41280;
  tmp_ivl_41288 <= y4(52);
  tmp_ivl_41289 <= new_AGEMA_signal_2386 & tmp_ivl_41288;
  LPM_q_ivl_41292 <= tmp_ivl_41294 & tmp_ivl_41289;
  tmp_ivl_41297 <= fresh(209);
  LPM_q_ivl_41299 <= tmp_ivl_41301 & tmp_ivl_41297;
  new_AGEMA_signal_3192 <= tmp_ivl_41305(1);
  tmp_ivl_41303 <= tmp_ivl_41305(0);
  tmp_ivl_41305 <= LPM_d0_ivl_41309(0 + 1 downto 0);
  tmp_ivl_41310 <= new_AGEMA_signal_2877 & SboxInst_n344;
  LPM_q_ivl_41313 <= tmp_ivl_41315 & tmp_ivl_41310;
  tmp_ivl_41318 <= y4(46);
  tmp_ivl_41319 <= new_AGEMA_signal_2407 & tmp_ivl_41318;
  LPM_q_ivl_41322 <= tmp_ivl_41324 & tmp_ivl_41319;
  tmp_ivl_41327 <= fresh(210);
  LPM_q_ivl_41329 <= tmp_ivl_41331 & tmp_ivl_41327;
  new_AGEMA_signal_3193 <= tmp_ivl_41335(1);
  tmp_ivl_41333 <= tmp_ivl_41335(0);
  tmp_ivl_41335 <= LPM_d0_ivl_41339(0 + 1 downto 0);
  tmp_ivl_41340 <= new_AGEMA_signal_2878 & SboxInst_n338;
  LPM_q_ivl_41343 <= tmp_ivl_41345 & tmp_ivl_41340;
  tmp_ivl_41348 <= y4(51);
  tmp_ivl_41349 <= new_AGEMA_signal_2389 & tmp_ivl_41348;
  LPM_q_ivl_41352 <= tmp_ivl_41354 & tmp_ivl_41349;
  tmp_ivl_41357 <= fresh(211);
  LPM_q_ivl_41359 <= tmp_ivl_41361 & tmp_ivl_41357;
  new_AGEMA_signal_3194 <= tmp_ivl_41365(1);
  tmp_ivl_41363 <= tmp_ivl_41365(0);
  tmp_ivl_41365 <= LPM_d0_ivl_41369(0 + 1 downto 0);
  tmp_ivl_41370 <= new_AGEMA_signal_2879 & SboxInst_n339;
  LPM_q_ivl_41373 <= tmp_ivl_41375 & tmp_ivl_41370;
  tmp_ivl_41378 <= y4(50);
  tmp_ivl_41379 <= new_AGEMA_signal_2392 & tmp_ivl_41378;
  LPM_q_ivl_41382 <= tmp_ivl_41384 & tmp_ivl_41379;
  tmp_ivl_41387 <= fresh(212);
  LPM_q_ivl_41389 <= tmp_ivl_41391 & tmp_ivl_41387;
  new_AGEMA_signal_3195 <= tmp_ivl_41395(1);
  tmp_ivl_41393 <= tmp_ivl_41395(0);
  tmp_ivl_41395 <= LPM_d0_ivl_41399(0 + 1 downto 0);
  tmp_ivl_41400 <= new_AGEMA_signal_2880 & SboxInst_n341;
  LPM_q_ivl_41403 <= tmp_ivl_41405 & tmp_ivl_41400;
  tmp_ivl_41408 <= y4(49);
  tmp_ivl_41409 <= new_AGEMA_signal_2398 & tmp_ivl_41408;
  LPM_q_ivl_41412 <= tmp_ivl_41414 & tmp_ivl_41409;
  tmp_ivl_41417 <= fresh(213);
  LPM_q_ivl_41419 <= tmp_ivl_41421 & tmp_ivl_41417;
  new_AGEMA_signal_3196 <= tmp_ivl_41425(1);
  tmp_ivl_41423 <= tmp_ivl_41425(0);
  tmp_ivl_41425 <= LPM_d0_ivl_41429(0 + 1 downto 0);
  tmp_ivl_41430 <= new_AGEMA_signal_2881 & SboxInst_n334;
  LPM_q_ivl_41433 <= tmp_ivl_41435 & tmp_ivl_41430;
  tmp_ivl_41438 <= y4(55);
  tmp_ivl_41439 <= new_AGEMA_signal_2377 & tmp_ivl_41438;
  LPM_q_ivl_41442 <= tmp_ivl_41444 & tmp_ivl_41439;
  tmp_ivl_41447 <= fresh(214);
  LPM_q_ivl_41449 <= tmp_ivl_41451 & tmp_ivl_41447;
  new_AGEMA_signal_3197 <= tmp_ivl_41455(1);
  tmp_ivl_41453 <= tmp_ivl_41455(0);
  tmp_ivl_41455 <= LPM_d0_ivl_41459(0 + 1 downto 0);
  tmp_ivl_41460 <= new_AGEMA_signal_2882 & SboxInst_n327;
  LPM_q_ivl_41463 <= tmp_ivl_41465 & tmp_ivl_41460;
  tmp_ivl_41468 <= y4(61);
  tmp_ivl_41469 <= new_AGEMA_signal_2356 & tmp_ivl_41468;
  LPM_q_ivl_41472 <= tmp_ivl_41474 & tmp_ivl_41469;
  tmp_ivl_41477 <= fresh(215);
  LPM_q_ivl_41479 <= tmp_ivl_41481 & tmp_ivl_41477;
  new_AGEMA_signal_3198 <= tmp_ivl_41485(1);
  tmp_ivl_41483 <= tmp_ivl_41485(0);
  tmp_ivl_41485 <= LPM_d0_ivl_41489(0 + 1 downto 0);
  tmp_ivl_41490 <= new_AGEMA_signal_2883 & SboxInst_n333;
  LPM_q_ivl_41493 <= tmp_ivl_41495 & tmp_ivl_41490;
  tmp_ivl_41498 <= y4(56);
  tmp_ivl_41499 <= new_AGEMA_signal_2374 & tmp_ivl_41498;
  LPM_q_ivl_41502 <= tmp_ivl_41504 & tmp_ivl_41499;
  tmp_ivl_41507 <= fresh(216);
  LPM_q_ivl_41509 <= tmp_ivl_41511 & tmp_ivl_41507;
  new_AGEMA_signal_3199 <= tmp_ivl_41515(1);
  tmp_ivl_41513 <= tmp_ivl_41515(0);
  tmp_ivl_41515 <= LPM_d0_ivl_41519(0 + 1 downto 0);
  tmp_ivl_41520 <= new_AGEMA_signal_2884 & SboxInst_n335;
  LPM_q_ivl_41523 <= tmp_ivl_41525 & tmp_ivl_41520;
  tmp_ivl_41528 <= y4(54);
  tmp_ivl_41529 <= new_AGEMA_signal_2380 & tmp_ivl_41528;
  LPM_q_ivl_41532 <= tmp_ivl_41534 & tmp_ivl_41529;
  tmp_ivl_41537 <= fresh(217);
  LPM_q_ivl_41539 <= tmp_ivl_41541 & tmp_ivl_41537;
  new_AGEMA_signal_3200 <= tmp_ivl_41545(1);
  tmp_ivl_41543 <= tmp_ivl_41545(0);
  tmp_ivl_41545 <= LPM_d0_ivl_41549(0 + 1 downto 0);
  tmp_ivl_41550 <= new_AGEMA_signal_2885 & SboxInst_n328;
  LPM_q_ivl_41553 <= tmp_ivl_41555 & tmp_ivl_41550;
  tmp_ivl_41558 <= y4(60);
  tmp_ivl_41559 <= new_AGEMA_signal_2359 & tmp_ivl_41558;
  LPM_q_ivl_41562 <= tmp_ivl_41564 & tmp_ivl_41559;
  tmp_ivl_41567 <= fresh(218);
  LPM_q_ivl_41569 <= tmp_ivl_41571 & tmp_ivl_41567;
  new_AGEMA_signal_3201 <= tmp_ivl_41575(1);
  tmp_ivl_41573 <= tmp_ivl_41575(0);
  tmp_ivl_41575 <= LPM_d0_ivl_41579(0 + 1 downto 0);
  tmp_ivl_41580 <= new_AGEMA_signal_2886 & SboxInst_n330;
  LPM_q_ivl_41583 <= tmp_ivl_41585 & tmp_ivl_41580;
  tmp_ivl_41588 <= y4(59);
  tmp_ivl_41589 <= new_AGEMA_signal_2365 & tmp_ivl_41588;
  LPM_q_ivl_41592 <= tmp_ivl_41594 & tmp_ivl_41589;
  tmp_ivl_41597 <= fresh(219);
  LPM_q_ivl_41599 <= tmp_ivl_41601 & tmp_ivl_41597;
  new_AGEMA_signal_3202 <= tmp_ivl_41605(1);
  tmp_ivl_41603 <= tmp_ivl_41605(0);
  tmp_ivl_41605 <= LPM_d0_ivl_41609(0 + 1 downto 0);
  tmp_ivl_41610 <= new_AGEMA_signal_2887 & SboxInst_n331;
  LPM_q_ivl_41613 <= tmp_ivl_41615 & tmp_ivl_41610;
  tmp_ivl_41618 <= y4(58);
  tmp_ivl_41619 <= new_AGEMA_signal_2368 & tmp_ivl_41618;
  LPM_q_ivl_41622 <= tmp_ivl_41624 & tmp_ivl_41619;
  tmp_ivl_41627 <= fresh(220);
  LPM_q_ivl_41629 <= tmp_ivl_41631 & tmp_ivl_41627;
  new_AGEMA_signal_3203 <= tmp_ivl_41635(1);
  tmp_ivl_41633 <= tmp_ivl_41635(0);
  tmp_ivl_41635 <= LPM_d0_ivl_41639(0 + 1 downto 0);
  tmp_ivl_41640 <= new_AGEMA_signal_2888 & SboxInst_n332;
  LPM_q_ivl_41643 <= tmp_ivl_41645 & tmp_ivl_41640;
  tmp_ivl_41648 <= y4(57);
  tmp_ivl_41649 <= new_AGEMA_signal_2371 & tmp_ivl_41648;
  LPM_q_ivl_41652 <= tmp_ivl_41654 & tmp_ivl_41649;
  tmp_ivl_41657 <= fresh(221);
  LPM_q_ivl_41659 <= tmp_ivl_41661 & tmp_ivl_41657;
  new_AGEMA_signal_3204 <= tmp_ivl_41665(1);
  tmp_ivl_41663 <= tmp_ivl_41665(0);
  tmp_ivl_41665 <= LPM_d0_ivl_41669(0 + 1 downto 0);
  tmp_ivl_41670 <= new_AGEMA_signal_2889 & SboxInst_n325;
  LPM_q_ivl_41673 <= tmp_ivl_41675 & tmp_ivl_41670;
  tmp_ivl_41678 <= y4(63);
  tmp_ivl_41679 <= new_AGEMA_signal_2350 & tmp_ivl_41678;
  LPM_q_ivl_41682 <= tmp_ivl_41684 & tmp_ivl_41679;
  tmp_ivl_41687 <= fresh(222);
  LPM_q_ivl_41689 <= tmp_ivl_41691 & tmp_ivl_41687;
  new_AGEMA_signal_3205 <= tmp_ivl_41695(1);
  tmp_ivl_41693 <= tmp_ivl_41695(0);
  tmp_ivl_41695 <= LPM_d0_ivl_41699(0 + 1 downto 0);
  tmp_ivl_41700 <= new_AGEMA_signal_2890 & SboxInst_n384;
  LPM_q_ivl_41703 <= tmp_ivl_41705 & tmp_ivl_41700;
  tmp_ivl_41708 <= y4(0);
  tmp_ivl_41709 <= new_AGEMA_signal_2527 & tmp_ivl_41708;
  LPM_q_ivl_41712 <= tmp_ivl_41714 & tmp_ivl_41709;
  tmp_ivl_41717 <= fresh(223);
  LPM_q_ivl_41719 <= tmp_ivl_41721 & tmp_ivl_41717;
  new_AGEMA_signal_3206 <= tmp_ivl_41725(1);
  tmp_ivl_41723 <= tmp_ivl_41725(0);
  tmp_ivl_41725 <= LPM_d0_ivl_41729(0 + 1 downto 0);
  tmp_ivl_41730 <= new_AGEMA_signal_2891 & SboxInst_n329;
  LPM_q_ivl_41733 <= tmp_ivl_41735 & tmp_ivl_41730;
  tmp_ivl_41738 <= y4(5);
  tmp_ivl_41739 <= new_AGEMA_signal_2362 & tmp_ivl_41738;
  LPM_q_ivl_41742 <= tmp_ivl_41744 & tmp_ivl_41739;
  tmp_ivl_41747 <= fresh(224);
  LPM_q_ivl_41749 <= tmp_ivl_41751 & tmp_ivl_41747;
  new_AGEMA_signal_3207 <= tmp_ivl_41755(1);
  tmp_ivl_41753 <= tmp_ivl_41755(0);
  tmp_ivl_41755 <= LPM_d0_ivl_41759(0 + 1 downto 0);
  tmp_ivl_41760 <= new_AGEMA_signal_2892 & SboxInst_n340;
  LPM_q_ivl_41763 <= tmp_ivl_41765 & tmp_ivl_41760;
  tmp_ivl_41768 <= y4(4);
  tmp_ivl_41769 <= new_AGEMA_signal_2395 & tmp_ivl_41768;
  LPM_q_ivl_41772 <= tmp_ivl_41774 & tmp_ivl_41769;
  tmp_ivl_41777 <= fresh(225);
  LPM_q_ivl_41779 <= tmp_ivl_41781 & tmp_ivl_41777;
  new_AGEMA_signal_3208 <= tmp_ivl_41785(1);
  tmp_ivl_41783 <= tmp_ivl_41785(0);
  tmp_ivl_41785 <= LPM_d0_ivl_41789(0 + 1 downto 0);
  tmp_ivl_41790 <= new_AGEMA_signal_2893 & SboxInst_n326;
  LPM_q_ivl_41793 <= tmp_ivl_41795 & tmp_ivl_41790;
  tmp_ivl_41798 <= y4(62);
  tmp_ivl_41799 <= new_AGEMA_signal_2353 & tmp_ivl_41798;
  LPM_q_ivl_41802 <= tmp_ivl_41804 & tmp_ivl_41799;
  tmp_ivl_41807 <= fresh(226);
  LPM_q_ivl_41809 <= tmp_ivl_41811 & tmp_ivl_41807;
  new_AGEMA_signal_3209 <= tmp_ivl_41815(1);
  tmp_ivl_41813 <= tmp_ivl_41815(0);
  tmp_ivl_41815 <= LPM_d0_ivl_41819(0 + 1 downto 0);
  tmp_ivl_41820 <= new_AGEMA_signal_2894 & SboxInst_n351;
  LPM_q_ivl_41823 <= tmp_ivl_41825 & tmp_ivl_41820;
  tmp_ivl_41828 <= y4(3);
  tmp_ivl_41829 <= new_AGEMA_signal_2428 & tmp_ivl_41828;
  LPM_q_ivl_41832 <= tmp_ivl_41834 & tmp_ivl_41829;
  tmp_ivl_41837 <= fresh(227);
  LPM_q_ivl_41839 <= tmp_ivl_41841 & tmp_ivl_41837;
  new_AGEMA_signal_3210 <= tmp_ivl_41845(1);
  tmp_ivl_41843 <= tmp_ivl_41845(0);
  tmp_ivl_41845 <= LPM_d0_ivl_41849(0 + 1 downto 0);
  tmp_ivl_41850 <= new_AGEMA_signal_2895 & SboxInst_n362;
  LPM_q_ivl_41853 <= tmp_ivl_41855 & tmp_ivl_41850;
  tmp_ivl_41858 <= y4(2);
  tmp_ivl_41859 <= new_AGEMA_signal_2461 & tmp_ivl_41858;
  LPM_q_ivl_41862 <= tmp_ivl_41864 & tmp_ivl_41859;
  tmp_ivl_41867 <= fresh(228);
  LPM_q_ivl_41869 <= tmp_ivl_41871 & tmp_ivl_41867;
  new_AGEMA_signal_3211 <= tmp_ivl_41875(1);
  tmp_ivl_41873 <= tmp_ivl_41875(0);
  tmp_ivl_41875 <= LPM_d0_ivl_41879(0 + 1 downto 0);
  tmp_ivl_41880 <= new_AGEMA_signal_2896 & SboxInst_n373;
  LPM_q_ivl_41883 <= tmp_ivl_41885 & tmp_ivl_41880;
  tmp_ivl_41888 <= y4(1);
  tmp_ivl_41889 <= new_AGEMA_signal_2494 & tmp_ivl_41888;
  LPM_q_ivl_41892 <= tmp_ivl_41894 & tmp_ivl_41889;
  tmp_ivl_41897 <= fresh(229);
  LPM_q_ivl_41899 <= tmp_ivl_41901 & tmp_ivl_41897;
  new_AGEMA_signal_3212 <= tmp_ivl_41905(1);
  tmp_ivl_41903 <= tmp_ivl_41905(0);
  tmp_ivl_41905 <= LPM_d0_ivl_41909(0 + 1 downto 0);
  tmp_ivl_41910 <= new_AGEMA_signal_2793 & n3253;
  LPM_q_ivl_41913 <= tmp_ivl_41915 & tmp_ivl_41910;
  tmp_ivl_41917 <= new_AGEMA_signal_2897 & SboxInst_n216;
  LPM_q_ivl_41920 <= tmp_ivl_41922 & tmp_ivl_41917;
  tmp_ivl_41925 <= fresh(230);
  LPM_q_ivl_41927 <= tmp_ivl_41929 & tmp_ivl_41925;
  new_AGEMA_signal_3213 <= tmp_ivl_41933(1);
  tmp_ivl_41931 <= tmp_ivl_41933(0);
  tmp_ivl_41933 <= LPM_d0_ivl_41937(0 + 1 downto 0);
  tmp_ivl_41938 <= new_AGEMA_signal_4433 & n3239;
  LPM_q_ivl_41941 <= tmp_ivl_41943 & tmp_ivl_41938;
  tmp_ivl_41945 <= new_AGEMA_signal_2899 & SboxInst_n195;
  LPM_q_ivl_41948 <= tmp_ivl_41950 & tmp_ivl_41945;
  tmp_ivl_41953 <= fresh(231);
  LPM_q_ivl_41955 <= tmp_ivl_41957 & tmp_ivl_41953;
  new_AGEMA_signal_4579 <= tmp_ivl_41961(1);
  tmp_ivl_41959 <= tmp_ivl_41961(0);
  tmp_ivl_41961 <= LPM_d0_ivl_41965(0 + 1 downto 0);
  tmp_ivl_41966 <= new_AGEMA_signal_2990 & n3232;
  LPM_q_ivl_41969 <= tmp_ivl_41971 & tmp_ivl_41966;
  tmp_ivl_41973 <= new_AGEMA_signal_2900 & SboxInst_n212;
  LPM_q_ivl_41976 <= tmp_ivl_41978 & tmp_ivl_41973;
  tmp_ivl_41981 <= fresh(232);
  LPM_q_ivl_41983 <= tmp_ivl_41985 & tmp_ivl_41981;
  new_AGEMA_signal_3583 <= tmp_ivl_41989(1);
  tmp_ivl_41987 <= tmp_ivl_41989(0);
  tmp_ivl_41989 <= LPM_d0_ivl_41993(0 + 1 downto 0);
  tmp_ivl_41994 <= new_AGEMA_signal_3826 & n3230;
  LPM_q_ivl_41997 <= tmp_ivl_41999 & tmp_ivl_41994;
  tmp_ivl_42001 <= new_AGEMA_signal_2901 & SboxInst_n196;
  LPM_q_ivl_42004 <= tmp_ivl_42006 & tmp_ivl_42001;
  tmp_ivl_42009 <= fresh(233);
  LPM_q_ivl_42011 <= tmp_ivl_42013 & tmp_ivl_42009;
  new_AGEMA_signal_4202 <= tmp_ivl_42017(1);
  tmp_ivl_42015 <= tmp_ivl_42017(0);
  tmp_ivl_42017 <= LPM_d0_ivl_42021(0 + 1 downto 0);
  tmp_ivl_42022 <= new_AGEMA_signal_2790 & n3254;
  LPM_q_ivl_42025 <= tmp_ivl_42027 & tmp_ivl_42022;
  tmp_ivl_42029 <= new_AGEMA_signal_2902 & SboxInst_n217;
  LPM_q_ivl_42032 <= tmp_ivl_42034 & tmp_ivl_42029;
  tmp_ivl_42037 <= fresh(234);
  LPM_q_ivl_42039 <= tmp_ivl_42041 & tmp_ivl_42037;
  new_AGEMA_signal_3214 <= tmp_ivl_42045(1);
  tmp_ivl_42043 <= tmp_ivl_42045(0);
  tmp_ivl_42045 <= LPM_d0_ivl_42049(0 + 1 downto 0);
  tmp_ivl_42050 <= new_AGEMA_signal_4432 & n3233;
  LPM_q_ivl_42053 <= tmp_ivl_42055 & tmp_ivl_42050;
  tmp_ivl_42057 <= new_AGEMA_signal_2904 & SboxInst_n223;
  LPM_q_ivl_42060 <= tmp_ivl_42062 & tmp_ivl_42057;
  tmp_ivl_42065 <= fresh(235);
  LPM_q_ivl_42067 <= tmp_ivl_42069 & tmp_ivl_42065;
  new_AGEMA_signal_4580 <= tmp_ivl_42073(1);
  tmp_ivl_42071 <= tmp_ivl_42073(0);
  tmp_ivl_42073 <= LPM_d0_ivl_42077(0 + 1 downto 0);
  tmp_ivl_42078 <= new_AGEMA_signal_2788 & n3255;
  LPM_q_ivl_42081 <= tmp_ivl_42083 & tmp_ivl_42078;
  tmp_ivl_42085 <= new_AGEMA_signal_2905 & SboxInst_n218;
  LPM_q_ivl_42088 <= tmp_ivl_42090 & tmp_ivl_42085;
  tmp_ivl_42093 <= fresh(236);
  LPM_q_ivl_42095 <= tmp_ivl_42097 & tmp_ivl_42093;
  new_AGEMA_signal_3215 <= tmp_ivl_42101(1);
  tmp_ivl_42099 <= tmp_ivl_42101(0);
  tmp_ivl_42101 <= LPM_d0_ivl_42105(0 + 1 downto 0);
  tmp_ivl_42106 <= new_AGEMA_signal_3824 & n3287;
  LPM_q_ivl_42109 <= tmp_ivl_42111 & tmp_ivl_42106;
  tmp_ivl_42113 <= new_AGEMA_signal_2906 & SboxInst_n234;
  LPM_q_ivl_42116 <= tmp_ivl_42118 & tmp_ivl_42113;
  tmp_ivl_42121 <= fresh(237);
  LPM_q_ivl_42123 <= tmp_ivl_42125 & tmp_ivl_42121;
  new_AGEMA_signal_4203 <= tmp_ivl_42129(1);
  tmp_ivl_42127 <= tmp_ivl_42129(0);
  tmp_ivl_42129 <= LPM_d0_ivl_42133(0 + 1 downto 0);
  tmp_ivl_42134 <= new_AGEMA_signal_3515 & n3231;
  LPM_q_ivl_42137 <= tmp_ivl_42139 & tmp_ivl_42134;
  tmp_ivl_42141 <= new_AGEMA_signal_2907 & SboxInst_n201;
  LPM_q_ivl_42144 <= tmp_ivl_42146 & tmp_ivl_42141;
  tmp_ivl_42149 <= fresh(238);
  LPM_q_ivl_42151 <= tmp_ivl_42153 & tmp_ivl_42149;
  new_AGEMA_signal_3889 <= tmp_ivl_42157(1);
  tmp_ivl_42155 <= tmp_ivl_42157(0);
  tmp_ivl_42157 <= LPM_d0_ivl_42161(0 + 1 downto 0);
  tmp_ivl_42162 <= new_AGEMA_signal_2786 & n3256;
  LPM_q_ivl_42165 <= tmp_ivl_42167 & tmp_ivl_42162;
  tmp_ivl_42169 <= new_AGEMA_signal_2908 & SboxInst_n219;
  LPM_q_ivl_42172 <= tmp_ivl_42174 & tmp_ivl_42169;
  tmp_ivl_42177 <= fresh(239);
  LPM_q_ivl_42179 <= tmp_ivl_42181 & tmp_ivl_42177;
  new_AGEMA_signal_3216 <= tmp_ivl_42185(1);
  tmp_ivl_42183 <= tmp_ivl_42185(0);
  tmp_ivl_42185 <= LPM_d0_ivl_42189(0 + 1 downto 0);
  tmp_ivl_42191 <= y2(1);
  tmp_ivl_42192 <= new_AGEMA_signal_3513 & tmp_ivl_42191;
  LPM_q_ivl_42195 <= tmp_ivl_42197 & tmp_ivl_42192;
  tmp_ivl_42199 <= new_AGEMA_signal_2909 & SboxInst_n245;
  LPM_q_ivl_42202 <= tmp_ivl_42204 & tmp_ivl_42199;
  tmp_ivl_42207 <= fresh(240);
  LPM_q_ivl_42209 <= tmp_ivl_42211 & tmp_ivl_42207;
  new_AGEMA_signal_3890 <= tmp_ivl_42215(1);
  tmp_ivl_42213 <= tmp_ivl_42215(0);
  tmp_ivl_42215 <= LPM_d0_ivl_42219(0 + 1 downto 0);
  tmp_ivl_42220 <= new_AGEMA_signal_2783 & n3257;
  LPM_q_ivl_42223 <= tmp_ivl_42225 & tmp_ivl_42220;
  tmp_ivl_42227 <= new_AGEMA_signal_2910 & SboxInst_n220;
  LPM_q_ivl_42230 <= tmp_ivl_42232 & tmp_ivl_42227;
  tmp_ivl_42235 <= fresh(241);
  LPM_q_ivl_42237 <= tmp_ivl_42239 & tmp_ivl_42235;
  new_AGEMA_signal_3217 <= tmp_ivl_42243(1);
  tmp_ivl_42241 <= tmp_ivl_42243(0);
  tmp_ivl_42243 <= LPM_d0_ivl_42247(0 + 1 downto 0);
  tmp_ivl_42249 <= y2(0);
  tmp_ivl_42250 <= new_AGEMA_signal_2989 & tmp_ivl_42249;
  LPM_q_ivl_42253 <= tmp_ivl_42255 & tmp_ivl_42250;
  tmp_ivl_42257 <= new_AGEMA_signal_2911 & SboxInst_n256;
  LPM_q_ivl_42260 <= tmp_ivl_42262 & tmp_ivl_42257;
  tmp_ivl_42265 <= fresh(242);
  LPM_q_ivl_42267 <= tmp_ivl_42269 & tmp_ivl_42265;
  new_AGEMA_signal_3584 <= tmp_ivl_42273(1);
  tmp_ivl_42271 <= tmp_ivl_42273(0);
  tmp_ivl_42273 <= LPM_d0_ivl_42277(0 + 1 downto 0);
  tmp_ivl_42278 <= new_AGEMA_signal_2846 & n3234;
  LPM_q_ivl_42281 <= tmp_ivl_42283 & tmp_ivl_42278;
  tmp_ivl_42285 <= new_AGEMA_signal_2912 & SboxInst_n197;
  LPM_q_ivl_42288 <= tmp_ivl_42290 & tmp_ivl_42285;
  tmp_ivl_42293 <= fresh(243);
  LPM_q_ivl_42295 <= tmp_ivl_42297 & tmp_ivl_42293;
  new_AGEMA_signal_3218 <= tmp_ivl_42301(1);
  tmp_ivl_42299 <= tmp_ivl_42301(0);
  tmp_ivl_42301 <= LPM_d0_ivl_42305(0 + 1 downto 0);
  tmp_ivl_42306 <= new_AGEMA_signal_2780 & n3258;
  LPM_q_ivl_42309 <= tmp_ivl_42311 & tmp_ivl_42306;
  tmp_ivl_42313 <= new_AGEMA_signal_2913 & SboxInst_n221;
  LPM_q_ivl_42316 <= tmp_ivl_42318 & tmp_ivl_42313;
  tmp_ivl_42321 <= fresh(244);
  LPM_q_ivl_42323 <= tmp_ivl_42325 & tmp_ivl_42321;
  new_AGEMA_signal_3219 <= tmp_ivl_42329(1);
  tmp_ivl_42327 <= tmp_ivl_42329(0);
  tmp_ivl_42329 <= LPM_d0_ivl_42333(0 + 1 downto 0);
  tmp_ivl_42334 <= new_AGEMA_signal_2778 & n3259;
  LPM_q_ivl_42337 <= tmp_ivl_42339 & tmp_ivl_42334;
  tmp_ivl_42341 <= new_AGEMA_signal_2914 & SboxInst_n222;
  LPM_q_ivl_42344 <= tmp_ivl_42346 & tmp_ivl_42341;
  tmp_ivl_42349 <= fresh(245);
  LPM_q_ivl_42351 <= tmp_ivl_42353 & tmp_ivl_42349;
  new_AGEMA_signal_3220 <= tmp_ivl_42357(1);
  tmp_ivl_42355 <= tmp_ivl_42357(0);
  tmp_ivl_42357 <= LPM_d0_ivl_42361(0 + 1 downto 0);
  tmp_ivl_42362 <= new_AGEMA_signal_2840 & n3235;
  LPM_q_ivl_42365 <= tmp_ivl_42367 & tmp_ivl_42362;
  tmp_ivl_42369 <= new_AGEMA_signal_2915 & SboxInst_n198;
  LPM_q_ivl_42372 <= tmp_ivl_42374 & tmp_ivl_42369;
  tmp_ivl_42377 <= fresh(246);
  LPM_q_ivl_42379 <= tmp_ivl_42381 & tmp_ivl_42377;
  new_AGEMA_signal_3221 <= tmp_ivl_42385(1);
  tmp_ivl_42383 <= tmp_ivl_42385(0);
  tmp_ivl_42385 <= LPM_d0_ivl_42389(0 + 1 downto 0);
  tmp_ivl_42390 <= new_AGEMA_signal_2775 & n3260;
  LPM_q_ivl_42393 <= tmp_ivl_42395 & tmp_ivl_42390;
  tmp_ivl_42397 <= new_AGEMA_signal_2916 & SboxInst_n224;
  LPM_q_ivl_42400 <= tmp_ivl_42402 & tmp_ivl_42397;
  tmp_ivl_42405 <= fresh(247);
  LPM_q_ivl_42407 <= tmp_ivl_42409 & tmp_ivl_42405;
  new_AGEMA_signal_3222 <= tmp_ivl_42413(1);
  tmp_ivl_42411 <= tmp_ivl_42413(0);
  tmp_ivl_42413 <= LPM_d0_ivl_42417(0 + 1 downto 0);
  tmp_ivl_42418 <= new_AGEMA_signal_2837 & n3236;
  LPM_q_ivl_42421 <= tmp_ivl_42423 & tmp_ivl_42418;
  tmp_ivl_42425 <= new_AGEMA_signal_2917 & SboxInst_n199;
  LPM_q_ivl_42428 <= tmp_ivl_42430 & tmp_ivl_42425;
  tmp_ivl_42433 <= fresh(248);
  LPM_q_ivl_42435 <= tmp_ivl_42437 & tmp_ivl_42433;
  new_AGEMA_signal_3223 <= tmp_ivl_42441(1);
  tmp_ivl_42439 <= tmp_ivl_42441(0);
  tmp_ivl_42441 <= LPM_d0_ivl_42445(0 + 1 downto 0);
  tmp_ivl_42446 <= new_AGEMA_signal_2742 & n3284;
  LPM_q_ivl_42449 <= tmp_ivl_42451 & tmp_ivl_42446;
  tmp_ivl_42453 <= new_AGEMA_signal_2918 & SboxInst_n250;
  LPM_q_ivl_42456 <= tmp_ivl_42458 & tmp_ivl_42453;
  tmp_ivl_42461 <= fresh(249);
  LPM_q_ivl_42463 <= tmp_ivl_42465 & tmp_ivl_42461;
  new_AGEMA_signal_3224 <= tmp_ivl_42469(1);
  tmp_ivl_42467 <= tmp_ivl_42469(0);
  tmp_ivl_42469 <= LPM_d0_ivl_42473(0 + 1 downto 0);
  tmp_ivl_42474 <= new_AGEMA_signal_2717 & n3288;
  LPM_q_ivl_42477 <= tmp_ivl_42479 & tmp_ivl_42474;
  tmp_ivl_42481 <= new_AGEMA_signal_2919 & SboxInst_n253;
  LPM_q_ivl_42484 <= tmp_ivl_42486 & tmp_ivl_42481;
  tmp_ivl_42489 <= fresh(250);
  LPM_q_ivl_42491 <= tmp_ivl_42493 & tmp_ivl_42489;
  new_AGEMA_signal_3225 <= tmp_ivl_42497(1);
  tmp_ivl_42495 <= tmp_ivl_42497(0);
  tmp_ivl_42497 <= LPM_d0_ivl_42501(0 + 1 downto 0);
  tmp_ivl_42502 <= new_AGEMA_signal_2813 & n3245;
  LPM_q_ivl_42505 <= tmp_ivl_42507 & tmp_ivl_42502;
  tmp_ivl_42509 <= new_AGEMA_signal_2920 & SboxInst_n207;
  LPM_q_ivl_42512 <= tmp_ivl_42514 & tmp_ivl_42509;
  tmp_ivl_42517 <= fresh(251);
  LPM_q_ivl_42519 <= tmp_ivl_42521 & tmp_ivl_42517;
  new_AGEMA_signal_3226 <= tmp_ivl_42525(1);
  tmp_ivl_42523 <= tmp_ivl_42525(0);
  tmp_ivl_42525 <= LPM_d0_ivl_42529(0 + 1 downto 0);
  tmp_ivl_42530 <= new_AGEMA_signal_2709 & n3289;
  LPM_q_ivl_42533 <= tmp_ivl_42535 & tmp_ivl_42530;
  tmp_ivl_42537 <= new_AGEMA_signal_2921 & SboxInst_n254;
  LPM_q_ivl_42540 <= tmp_ivl_42542 & tmp_ivl_42537;
  tmp_ivl_42545 <= fresh(252);
  LPM_q_ivl_42547 <= tmp_ivl_42549 & tmp_ivl_42545;
  new_AGEMA_signal_3227 <= tmp_ivl_42553(1);
  tmp_ivl_42551 <= tmp_ivl_42553(0);
  tmp_ivl_42553 <= LPM_d0_ivl_42557(0 + 1 downto 0);
  tmp_ivl_42558 <= new_AGEMA_signal_2733 & n3285;
  LPM_q_ivl_42561 <= tmp_ivl_42563 & tmp_ivl_42558;
  tmp_ivl_42565 <= new_AGEMA_signal_2922 & SboxInst_n251;
  LPM_q_ivl_42568 <= tmp_ivl_42570 & tmp_ivl_42565;
  tmp_ivl_42573 <= fresh(253);
  LPM_q_ivl_42575 <= tmp_ivl_42577 & tmp_ivl_42573;
  new_AGEMA_signal_3228 <= tmp_ivl_42581(1);
  tmp_ivl_42579 <= tmp_ivl_42581(0);
  tmp_ivl_42581 <= LPM_d0_ivl_42585(0 + 1 downto 0);
  tmp_ivl_42586 <= new_AGEMA_signal_2810 & n3246;
  LPM_q_ivl_42589 <= tmp_ivl_42591 & tmp_ivl_42586;
  tmp_ivl_42593 <= new_AGEMA_signal_2923 & SboxInst_n208;
  LPM_q_ivl_42596 <= tmp_ivl_42598 & tmp_ivl_42593;
  tmp_ivl_42601 <= fresh(254);
  LPM_q_ivl_42603 <= tmp_ivl_42605 & tmp_ivl_42601;
  new_AGEMA_signal_3229 <= tmp_ivl_42609(1);
  tmp_ivl_42607 <= tmp_ivl_42609(0);
  tmp_ivl_42609 <= LPM_d0_ivl_42613(0 + 1 downto 0);
  tmp_ivl_42614 <= new_AGEMA_signal_2704 & n3290;
  LPM_q_ivl_42617 <= tmp_ivl_42619 & tmp_ivl_42614;
  tmp_ivl_42621 <= new_AGEMA_signal_2924 & SboxInst_n255;
  LPM_q_ivl_42624 <= tmp_ivl_42626 & tmp_ivl_42621;
  tmp_ivl_42629 <= fresh(255);
  LPM_q_ivl_42631 <= tmp_ivl_42633 & tmp_ivl_42629;
  new_AGEMA_signal_3230 <= tmp_ivl_42637(1);
  tmp_ivl_42635 <= tmp_ivl_42637(0);
  tmp_ivl_42637 <= LPM_d0_ivl_42641(0 + 1 downto 0);
  tmp_ivl_42642 <= new_AGEMA_signal_2727 & n3286;
  LPM_q_ivl_42645 <= tmp_ivl_42647 & tmp_ivl_42642;
  tmp_ivl_42649 <= new_AGEMA_signal_2925 & SboxInst_n252;
  LPM_q_ivl_42652 <= tmp_ivl_42654 & tmp_ivl_42649;
  tmp_ivl_42657 <= fresh(256);
  LPM_q_ivl_42659 <= tmp_ivl_42661 & tmp_ivl_42657;
  new_AGEMA_signal_3231 <= tmp_ivl_42665(1);
  tmp_ivl_42663 <= tmp_ivl_42665(0);
  tmp_ivl_42665 <= LPM_d0_ivl_42669(0 + 1 downto 0);
  tmp_ivl_42670 <= new_AGEMA_signal_2807 & n3247;
  LPM_q_ivl_42673 <= tmp_ivl_42675 & tmp_ivl_42670;
  tmp_ivl_42677 <= new_AGEMA_signal_2926 & SboxInst_n209;
  LPM_q_ivl_42680 <= tmp_ivl_42682 & tmp_ivl_42677;
  tmp_ivl_42685 <= fresh(257);
  LPM_q_ivl_42687 <= tmp_ivl_42689 & tmp_ivl_42685;
  new_AGEMA_signal_3232 <= tmp_ivl_42693(1);
  tmp_ivl_42691 <= tmp_ivl_42693(0);
  tmp_ivl_42693 <= LPM_d0_ivl_42697(0 + 1 downto 0);
  tmp_ivl_42698 <= new_AGEMA_signal_2692 & n3291;
  LPM_q_ivl_42701 <= tmp_ivl_42703 & tmp_ivl_42698;
  tmp_ivl_42705 <= new_AGEMA_signal_2927 & SboxInst_n193;
  LPM_q_ivl_42708 <= tmp_ivl_42710 & tmp_ivl_42705;
  tmp_ivl_42713 <= fresh(258);
  LPM_q_ivl_42715 <= tmp_ivl_42717 & tmp_ivl_42713;
  new_AGEMA_signal_3233 <= tmp_ivl_42721(1);
  tmp_ivl_42719 <= tmp_ivl_42721(0);
  tmp_ivl_42721 <= LPM_d0_ivl_42725(0 + 1 downto 0);
  tmp_ivl_42726 <= new_AGEMA_signal_2805 & n3248;
  LPM_q_ivl_42729 <= tmp_ivl_42731 & tmp_ivl_42726;
  tmp_ivl_42733 <= new_AGEMA_signal_2928 & SboxInst_n210;
  LPM_q_ivl_42736 <= tmp_ivl_42738 & tmp_ivl_42733;
  tmp_ivl_42741 <= fresh(259);
  LPM_q_ivl_42743 <= tmp_ivl_42745 & tmp_ivl_42741;
  new_AGEMA_signal_3234 <= tmp_ivl_42749(1);
  tmp_ivl_42747 <= tmp_ivl_42749(0);
  tmp_ivl_42749 <= LPM_d0_ivl_42753(0 + 1 downto 0);
  tmp_ivl_42754 <= new_AGEMA_signal_2834 & n3237;
  LPM_q_ivl_42757 <= tmp_ivl_42759 & tmp_ivl_42754;
  tmp_ivl_42761 <= new_AGEMA_signal_2929 & SboxInst_n194;
  LPM_q_ivl_42764 <= tmp_ivl_42766 & tmp_ivl_42761;
  tmp_ivl_42769 <= fresh(260);
  LPM_q_ivl_42771 <= tmp_ivl_42773 & tmp_ivl_42769;
  new_AGEMA_signal_3235 <= tmp_ivl_42777(1);
  tmp_ivl_42775 <= tmp_ivl_42777(0);
  tmp_ivl_42777 <= LPM_d0_ivl_42781(0 + 1 downto 0);
  tmp_ivl_42782 <= new_AGEMA_signal_2803 & n3249;
  LPM_q_ivl_42785 <= tmp_ivl_42787 & tmp_ivl_42782;
  tmp_ivl_42789 <= new_AGEMA_signal_2930 & SboxInst_n211;
  LPM_q_ivl_42792 <= tmp_ivl_42794 & tmp_ivl_42789;
  tmp_ivl_42797 <= fresh(261);
  LPM_q_ivl_42799 <= tmp_ivl_42801 & tmp_ivl_42797;
  new_AGEMA_signal_3236 <= tmp_ivl_42805(1);
  tmp_ivl_42803 <= tmp_ivl_42805(0);
  tmp_ivl_42805 <= LPM_d0_ivl_42809(0 + 1 downto 0);
  tmp_ivl_42810 <= new_AGEMA_signal_2800 & n3250;
  LPM_q_ivl_42813 <= tmp_ivl_42815 & tmp_ivl_42810;
  tmp_ivl_42817 <= new_AGEMA_signal_2931 & SboxInst_n213;
  LPM_q_ivl_42820 <= tmp_ivl_42822 & tmp_ivl_42817;
  tmp_ivl_42825 <= fresh(262);
  LPM_q_ivl_42827 <= tmp_ivl_42829 & tmp_ivl_42825;
  new_AGEMA_signal_3237 <= tmp_ivl_42833(1);
  tmp_ivl_42831 <= tmp_ivl_42833(0);
  tmp_ivl_42833 <= LPM_d0_ivl_42837(0 + 1 downto 0);
  tmp_ivl_42838 <= new_AGEMA_signal_2797 & n3251;
  LPM_q_ivl_42841 <= tmp_ivl_42843 & tmp_ivl_42838;
  tmp_ivl_42845 <= new_AGEMA_signal_2932 & SboxInst_n214;
  LPM_q_ivl_42848 <= tmp_ivl_42850 & tmp_ivl_42845;
  tmp_ivl_42853 <= fresh(263);
  LPM_q_ivl_42855 <= tmp_ivl_42857 & tmp_ivl_42853;
  new_AGEMA_signal_3238 <= tmp_ivl_42861(1);
  tmp_ivl_42859 <= tmp_ivl_42861(0);
  tmp_ivl_42861 <= LPM_d0_ivl_42865(0 + 1 downto 0);
  tmp_ivl_42866 <= new_AGEMA_signal_2795 & n3252;
  LPM_q_ivl_42869 <= tmp_ivl_42871 & tmp_ivl_42866;
  tmp_ivl_42873 <= new_AGEMA_signal_2933 & SboxInst_n215;
  LPM_q_ivl_42876 <= tmp_ivl_42878 & tmp_ivl_42873;
  tmp_ivl_42881 <= fresh(264);
  LPM_q_ivl_42883 <= tmp_ivl_42885 & tmp_ivl_42881;
  new_AGEMA_signal_3239 <= tmp_ivl_42889(1);
  tmp_ivl_42887 <= tmp_ivl_42889(0);
  tmp_ivl_42889 <= LPM_d0_ivl_42893(0 + 1 downto 0);
  tmp_ivl_42894 <= new_AGEMA_signal_2701 & n3279;
  LPM_q_ivl_42897 <= tmp_ivl_42899 & tmp_ivl_42894;
  tmp_ivl_42901 <= new_AGEMA_signal_2934 & SboxInst_n244;
  LPM_q_ivl_42904 <= tmp_ivl_42906 & tmp_ivl_42901;
  tmp_ivl_42909 <= fresh(265);
  LPM_q_ivl_42911 <= tmp_ivl_42913 & tmp_ivl_42909;
  new_AGEMA_signal_3240 <= tmp_ivl_42917(1);
  tmp_ivl_42915 <= tmp_ivl_42917(0);
  tmp_ivl_42917 <= LPM_d0_ivl_42921(0 + 1 downto 0);
  tmp_ivl_42922 <= new_AGEMA_signal_2724 & n3276;
  LPM_q_ivl_42925 <= tmp_ivl_42927 & tmp_ivl_42922;
  tmp_ivl_42929 <= new_AGEMA_signal_2935 & SboxInst_n241;
  LPM_q_ivl_42932 <= tmp_ivl_42934 & tmp_ivl_42929;
  tmp_ivl_42937 <= fresh(266);
  LPM_q_ivl_42939 <= tmp_ivl_42941 & tmp_ivl_42937;
  new_AGEMA_signal_3241 <= tmp_ivl_42945(1);
  tmp_ivl_42943 <= tmp_ivl_42945(0);
  tmp_ivl_42945 <= LPM_d0_ivl_42949(0 + 1 downto 0);
  tmp_ivl_42950 <= new_AGEMA_signal_2695 & n3280;
  LPM_q_ivl_42953 <= tmp_ivl_42955 & tmp_ivl_42950;
  tmp_ivl_42957 <= new_AGEMA_signal_2936 & SboxInst_n246;
  LPM_q_ivl_42960 <= tmp_ivl_42962 & tmp_ivl_42957;
  tmp_ivl_42965 <= fresh(267);
  LPM_q_ivl_42967 <= tmp_ivl_42969 & tmp_ivl_42965;
  new_AGEMA_signal_3242 <= tmp_ivl_42973(1);
  tmp_ivl_42971 <= tmp_ivl_42973(0);
  tmp_ivl_42973 <= LPM_d0_ivl_42977(0 + 1 downto 0);
  tmp_ivl_42978 <= new_AGEMA_signal_2719 & n3277;
  LPM_q_ivl_42981 <= tmp_ivl_42983 & tmp_ivl_42978;
  tmp_ivl_42985 <= new_AGEMA_signal_2937 & SboxInst_n242;
  LPM_q_ivl_42988 <= tmp_ivl_42990 & tmp_ivl_42985;
  tmp_ivl_42993 <= fresh(268);
  LPM_q_ivl_42995 <= tmp_ivl_42997 & tmp_ivl_42993;
  new_AGEMA_signal_3243 <= tmp_ivl_43001(1);
  tmp_ivl_42999 <= tmp_ivl_43001(0);
  tmp_ivl_43001 <= LPM_d0_ivl_43005(0 + 1 downto 0);
  tmp_ivl_43006 <= new_AGEMA_signal_2828 & n3238;
  LPM_q_ivl_43009 <= tmp_ivl_43011 & tmp_ivl_43006;
  tmp_ivl_43013 <= new_AGEMA_signal_2938 & SboxInst_n200;
  LPM_q_ivl_43016 <= tmp_ivl_43018 & tmp_ivl_43013;
  tmp_ivl_43021 <= fresh(269);
  LPM_q_ivl_43023 <= tmp_ivl_43025 & tmp_ivl_43021;
  new_AGEMA_signal_3244 <= tmp_ivl_43029(1);
  tmp_ivl_43027 <= tmp_ivl_43029(0);
  tmp_ivl_43029 <= LPM_d0_ivl_43033(0 + 1 downto 0);
  tmp_ivl_43034 <= new_AGEMA_signal_2712 & n3278;
  LPM_q_ivl_43037 <= tmp_ivl_43039 & tmp_ivl_43034;
  tmp_ivl_43041 <= new_AGEMA_signal_2939 & SboxInst_n243;
  LPM_q_ivl_43044 <= tmp_ivl_43046 & tmp_ivl_43041;
  tmp_ivl_43049 <= fresh(270);
  LPM_q_ivl_43051 <= tmp_ivl_43053 & tmp_ivl_43049;
  new_AGEMA_signal_3245 <= tmp_ivl_43057(1);
  tmp_ivl_43055 <= tmp_ivl_43057(0);
  tmp_ivl_43057 <= LPM_d0_ivl_43061(0 + 1 downto 0);
  tmp_ivl_43062 <= new_AGEMA_signal_2760 & n3281;
  LPM_q_ivl_43065 <= tmp_ivl_43067 & tmp_ivl_43062;
  tmp_ivl_43069 <= new_AGEMA_signal_2940 & SboxInst_n247;
  LPM_q_ivl_43072 <= tmp_ivl_43074 & tmp_ivl_43069;
  tmp_ivl_43077 <= fresh(271);
  LPM_q_ivl_43079 <= tmp_ivl_43081 & tmp_ivl_43077;
  new_AGEMA_signal_3246 <= tmp_ivl_43085(1);
  tmp_ivl_43083 <= tmp_ivl_43085(0);
  tmp_ivl_43085 <= LPM_d0_ivl_43089(0 + 1 downto 0);
  tmp_ivl_43090 <= new_AGEMA_signal_2825 & n3240;
  LPM_q_ivl_43093 <= tmp_ivl_43095 & tmp_ivl_43090;
  tmp_ivl_43097 <= new_AGEMA_signal_2941 & SboxInst_n202;
  LPM_q_ivl_43100 <= tmp_ivl_43102 & tmp_ivl_43097;
  tmp_ivl_43105 <= fresh(272);
  LPM_q_ivl_43107 <= tmp_ivl_43109 & tmp_ivl_43105;
  new_AGEMA_signal_3247 <= tmp_ivl_43113(1);
  tmp_ivl_43111 <= tmp_ivl_43113(0);
  tmp_ivl_43113 <= LPM_d0_ivl_43117(0 + 1 downto 0);
  tmp_ivl_43118 <= new_AGEMA_signal_2755 & n3282;
  LPM_q_ivl_43121 <= tmp_ivl_43123 & tmp_ivl_43118;
  tmp_ivl_43125 <= new_AGEMA_signal_2942 & SboxInst_n248;
  LPM_q_ivl_43128 <= tmp_ivl_43130 & tmp_ivl_43125;
  tmp_ivl_43133 <= fresh(273);
  LPM_q_ivl_43135 <= tmp_ivl_43137 & tmp_ivl_43133;
  new_AGEMA_signal_3248 <= tmp_ivl_43141(1);
  tmp_ivl_43139 <= tmp_ivl_43141(0);
  tmp_ivl_43141 <= LPM_d0_ivl_43145(0 + 1 downto 0);
  tmp_ivl_43146 <= new_AGEMA_signal_2823 & n3241;
  LPM_q_ivl_43149 <= tmp_ivl_43151 & tmp_ivl_43146;
  tmp_ivl_43153 <= new_AGEMA_signal_2943 & SboxInst_n203;
  LPM_q_ivl_43156 <= tmp_ivl_43158 & tmp_ivl_43153;
  tmp_ivl_43161 <= fresh(274);
  LPM_q_ivl_43163 <= tmp_ivl_43165 & tmp_ivl_43161;
  new_AGEMA_signal_3249 <= tmp_ivl_43169(1);
  tmp_ivl_43167 <= tmp_ivl_43169(0);
  tmp_ivl_43169 <= LPM_d0_ivl_43173(0 + 1 downto 0);
  tmp_ivl_43174 <= new_AGEMA_signal_2750 & n3283;
  LPM_q_ivl_43177 <= tmp_ivl_43179 & tmp_ivl_43174;
  tmp_ivl_43181 <= new_AGEMA_signal_2944 & SboxInst_n249;
  LPM_q_ivl_43184 <= tmp_ivl_43186 & tmp_ivl_43181;
  tmp_ivl_43189 <= fresh(275);
  LPM_q_ivl_43191 <= tmp_ivl_43193 & tmp_ivl_43189;
  new_AGEMA_signal_3250 <= tmp_ivl_43197(1);
  tmp_ivl_43195 <= tmp_ivl_43197(0);
  tmp_ivl_43197 <= LPM_d0_ivl_43201(0 + 1 downto 0);
  tmp_ivl_43202 <= new_AGEMA_signal_2821 & n3242;
  LPM_q_ivl_43205 <= tmp_ivl_43207 & tmp_ivl_43202;
  tmp_ivl_43209 <= new_AGEMA_signal_2945 & SboxInst_n204;
  LPM_q_ivl_43212 <= tmp_ivl_43214 & tmp_ivl_43209;
  tmp_ivl_43217 <= fresh(276);
  LPM_q_ivl_43219 <= tmp_ivl_43221 & tmp_ivl_43217;
  new_AGEMA_signal_3251 <= tmp_ivl_43225(1);
  tmp_ivl_43223 <= tmp_ivl_43225(0);
  tmp_ivl_43225 <= LPM_d0_ivl_43229(0 + 1 downto 0);
  tmp_ivl_43230 <= new_AGEMA_signal_2819 & n3243;
  LPM_q_ivl_43233 <= tmp_ivl_43235 & tmp_ivl_43230;
  tmp_ivl_43237 <= new_AGEMA_signal_2946 & SboxInst_n205;
  LPM_q_ivl_43240 <= tmp_ivl_43242 & tmp_ivl_43237;
  tmp_ivl_43245 <= fresh(277);
  LPM_q_ivl_43247 <= tmp_ivl_43249 & tmp_ivl_43245;
  new_AGEMA_signal_3252 <= tmp_ivl_43253(1);
  tmp_ivl_43251 <= tmp_ivl_43253(0);
  tmp_ivl_43253 <= LPM_d0_ivl_43257(0 + 1 downto 0);
  tmp_ivl_43258 <= new_AGEMA_signal_2816 & n3244;
  LPM_q_ivl_43261 <= tmp_ivl_43263 & tmp_ivl_43258;
  tmp_ivl_43265 <= new_AGEMA_signal_2947 & SboxInst_n206;
  LPM_q_ivl_43268 <= tmp_ivl_43270 & tmp_ivl_43265;
  tmp_ivl_43273 <= fresh(278);
  LPM_q_ivl_43275 <= tmp_ivl_43277 & tmp_ivl_43273;
  new_AGEMA_signal_3253 <= tmp_ivl_43281(1);
  tmp_ivl_43279 <= tmp_ivl_43281(0);
  tmp_ivl_43281 <= LPM_d0_ivl_43285(0 + 1 downto 0);
  tmp_ivl_43286 <= new_AGEMA_signal_2739 & n3268;
  LPM_q_ivl_43289 <= tmp_ivl_43291 & tmp_ivl_43286;
  tmp_ivl_43293 <= new_AGEMA_signal_2948 & SboxInst_n232;
  LPM_q_ivl_43296 <= tmp_ivl_43298 & tmp_ivl_43293;
  tmp_ivl_43301 <= fresh(279);
  LPM_q_ivl_43303 <= tmp_ivl_43305 & tmp_ivl_43301;
  new_AGEMA_signal_3254 <= tmp_ivl_43309(1);
  tmp_ivl_43307 <= tmp_ivl_43309(0);
  tmp_ivl_43309 <= LPM_d0_ivl_43313(0 + 1 downto 0);
  tmp_ivl_43314 <= new_AGEMA_signal_2714 & n3271;
  LPM_q_ivl_43317 <= tmp_ivl_43319 & tmp_ivl_43314;
  tmp_ivl_43321 <= new_AGEMA_signal_2949 & SboxInst_n236;
  LPM_q_ivl_43324 <= tmp_ivl_43326 & tmp_ivl_43321;
  tmp_ivl_43329 <= fresh(280);
  LPM_q_ivl_43331 <= tmp_ivl_43333 & tmp_ivl_43329;
  new_AGEMA_signal_3255 <= tmp_ivl_43337(1);
  tmp_ivl_43335 <= tmp_ivl_43337(0);
  tmp_ivl_43337 <= LPM_d0_ivl_43341(0 + 1 downto 0);
  tmp_ivl_43342 <= new_AGEMA_signal_2730 & n3269;
  LPM_q_ivl_43345 <= tmp_ivl_43347 & tmp_ivl_43342;
  tmp_ivl_43349 <= new_AGEMA_signal_2950 & SboxInst_n233;
  LPM_q_ivl_43352 <= tmp_ivl_43354 & tmp_ivl_43349;
  tmp_ivl_43357 <= fresh(281);
  LPM_q_ivl_43359 <= tmp_ivl_43361 & tmp_ivl_43357;
  new_AGEMA_signal_3256 <= tmp_ivl_43365(1);
  tmp_ivl_43363 <= tmp_ivl_43365(0);
  tmp_ivl_43365 <= LPM_d0_ivl_43369(0 + 1 downto 0);
  tmp_ivl_43370 <= new_AGEMA_signal_2707 & n3272;
  LPM_q_ivl_43373 <= tmp_ivl_43375 & tmp_ivl_43370;
  tmp_ivl_43377 <= new_AGEMA_signal_2951 & SboxInst_n237;
  LPM_q_ivl_43380 <= tmp_ivl_43382 & tmp_ivl_43377;
  tmp_ivl_43385 <= fresh(282);
  LPM_q_ivl_43387 <= tmp_ivl_43389 & tmp_ivl_43385;
  new_AGEMA_signal_3257 <= tmp_ivl_43393(1);
  tmp_ivl_43391 <= tmp_ivl_43393(0);
  tmp_ivl_43393 <= LPM_d0_ivl_43397(0 + 1 downto 0);
  tmp_ivl_43398 <= new_AGEMA_signal_2698 & n3273;
  LPM_q_ivl_43401 <= tmp_ivl_43403 & tmp_ivl_43398;
  tmp_ivl_43405 <= new_AGEMA_signal_2952 & SboxInst_n238;
  LPM_q_ivl_43408 <= tmp_ivl_43410 & tmp_ivl_43405;
  tmp_ivl_43413 <= fresh(283);
  LPM_q_ivl_43415 <= tmp_ivl_43417 & tmp_ivl_43413;
  new_AGEMA_signal_3258 <= tmp_ivl_43421(1);
  tmp_ivl_43419 <= tmp_ivl_43421(0);
  tmp_ivl_43421 <= LPM_d0_ivl_43425(0 + 1 downto 0);
  tmp_ivl_43426 <= new_AGEMA_signal_2721 & n3270;
  LPM_q_ivl_43429 <= tmp_ivl_43431 & tmp_ivl_43426;
  tmp_ivl_43433 <= new_AGEMA_signal_2953 & SboxInst_n235;
  LPM_q_ivl_43436 <= tmp_ivl_43438 & tmp_ivl_43433;
  tmp_ivl_43441 <= fresh(284);
  LPM_q_ivl_43443 <= tmp_ivl_43445 & tmp_ivl_43441;
  new_AGEMA_signal_3259 <= tmp_ivl_43449(1);
  tmp_ivl_43447 <= tmp_ivl_43449(0);
  tmp_ivl_43449 <= LPM_d0_ivl_43453(0 + 1 downto 0);
  tmp_ivl_43454 <= new_AGEMA_signal_2744 & n3274;
  LPM_q_ivl_43457 <= tmp_ivl_43459 & tmp_ivl_43454;
  tmp_ivl_43461 <= new_AGEMA_signal_2954 & SboxInst_n239;
  LPM_q_ivl_43464 <= tmp_ivl_43466 & tmp_ivl_43461;
  tmp_ivl_43469 <= fresh(285);
  LPM_q_ivl_43471 <= tmp_ivl_43473 & tmp_ivl_43469;
  new_AGEMA_signal_3260 <= tmp_ivl_43477(1);
  tmp_ivl_43475 <= tmp_ivl_43477(0);
  tmp_ivl_43477 <= LPM_d0_ivl_43481(0 + 1 downto 0);
  tmp_ivl_43482 <= new_AGEMA_signal_2736 & n3275;
  LPM_q_ivl_43485 <= tmp_ivl_43487 & tmp_ivl_43482;
  tmp_ivl_43489 <= new_AGEMA_signal_2955 & SboxInst_n240;
  LPM_q_ivl_43492 <= tmp_ivl_43494 & tmp_ivl_43489;
  tmp_ivl_43497 <= fresh(286);
  LPM_q_ivl_43499 <= tmp_ivl_43501 & tmp_ivl_43497;
  new_AGEMA_signal_3261 <= tmp_ivl_43505(1);
  tmp_ivl_43503 <= tmp_ivl_43505(0);
  tmp_ivl_43505 <= LPM_d0_ivl_43509(0 + 1 downto 0);
  tmp_ivl_43510 <= new_AGEMA_signal_2766 & n3263;
  LPM_q_ivl_43513 <= tmp_ivl_43515 & tmp_ivl_43510;
  tmp_ivl_43517 <= new_AGEMA_signal_2956 & SboxInst_n227;
  LPM_q_ivl_43520 <= tmp_ivl_43522 & tmp_ivl_43517;
  tmp_ivl_43525 <= fresh(287);
  LPM_q_ivl_43527 <= tmp_ivl_43529 & tmp_ivl_43525;
  new_AGEMA_signal_3262 <= tmp_ivl_43533(1);
  tmp_ivl_43531 <= tmp_ivl_43533(0);
  tmp_ivl_43533 <= LPM_d0_ivl_43537(0 + 1 downto 0);
  tmp_ivl_43538 <= new_AGEMA_signal_2763 & n3264;
  LPM_q_ivl_43541 <= tmp_ivl_43543 & tmp_ivl_43538;
  tmp_ivl_43545 <= new_AGEMA_signal_2957 & SboxInst_n228;
  LPM_q_ivl_43548 <= tmp_ivl_43550 & tmp_ivl_43545;
  tmp_ivl_43553 <= fresh(288);
  LPM_q_ivl_43555 <= tmp_ivl_43557 & tmp_ivl_43553;
  new_AGEMA_signal_3263 <= tmp_ivl_43561(1);
  tmp_ivl_43559 <= tmp_ivl_43561(0);
  tmp_ivl_43561 <= LPM_d0_ivl_43565(0 + 1 downto 0);
  tmp_ivl_43566 <= new_AGEMA_signal_2772 & n3261;
  LPM_q_ivl_43569 <= tmp_ivl_43571 & tmp_ivl_43566;
  tmp_ivl_43573 <= new_AGEMA_signal_2958 & SboxInst_n225;
  LPM_q_ivl_43576 <= tmp_ivl_43578 & tmp_ivl_43573;
  tmp_ivl_43581 <= fresh(289);
  LPM_q_ivl_43583 <= tmp_ivl_43585 & tmp_ivl_43581;
  new_AGEMA_signal_3264 <= tmp_ivl_43589(1);
  tmp_ivl_43587 <= tmp_ivl_43589(0);
  tmp_ivl_43589 <= LPM_d0_ivl_43593(0 + 1 downto 0);
  tmp_ivl_43594 <= new_AGEMA_signal_2758 & n3265;
  LPM_q_ivl_43597 <= tmp_ivl_43599 & tmp_ivl_43594;
  tmp_ivl_43601 <= new_AGEMA_signal_2959 & SboxInst_n229;
  LPM_q_ivl_43604 <= tmp_ivl_43606 & tmp_ivl_43601;
  tmp_ivl_43609 <= fresh(290);
  LPM_q_ivl_43611 <= tmp_ivl_43613 & tmp_ivl_43609;
  new_AGEMA_signal_3265 <= tmp_ivl_43617(1);
  tmp_ivl_43615 <= tmp_ivl_43617(0);
  tmp_ivl_43617 <= LPM_d0_ivl_43621(0 + 1 downto 0);
  tmp_ivl_43622 <= new_AGEMA_signal_2769 & n3262;
  LPM_q_ivl_43625 <= tmp_ivl_43627 & tmp_ivl_43622;
  tmp_ivl_43629 <= new_AGEMA_signal_2960 & SboxInst_n226;
  LPM_q_ivl_43632 <= tmp_ivl_43634 & tmp_ivl_43629;
  tmp_ivl_43637 <= fresh(291);
  LPM_q_ivl_43639 <= tmp_ivl_43641 & tmp_ivl_43637;
  new_AGEMA_signal_3266 <= tmp_ivl_43645(1);
  tmp_ivl_43643 <= tmp_ivl_43645(0);
  tmp_ivl_43645 <= LPM_d0_ivl_43649(0 + 1 downto 0);
  tmp_ivl_43650 <= new_AGEMA_signal_2753 & n3266;
  LPM_q_ivl_43653 <= tmp_ivl_43655 & tmp_ivl_43650;
  tmp_ivl_43657 <= new_AGEMA_signal_2961 & SboxInst_n230;
  LPM_q_ivl_43660 <= tmp_ivl_43662 & tmp_ivl_43657;
  tmp_ivl_43665 <= fresh(292);
  LPM_q_ivl_43667 <= tmp_ivl_43669 & tmp_ivl_43665;
  new_AGEMA_signal_3267 <= tmp_ivl_43673(1);
  tmp_ivl_43671 <= tmp_ivl_43673(0);
  tmp_ivl_43673 <= LPM_d0_ivl_43677(0 + 1 downto 0);
  tmp_ivl_43678 <= new_AGEMA_signal_2747 & n3267;
  LPM_q_ivl_43681 <= tmp_ivl_43683 & tmp_ivl_43678;
  tmp_ivl_43685 <= new_AGEMA_signal_2962 & SboxInst_n231;
  LPM_q_ivl_43688 <= tmp_ivl_43690 & tmp_ivl_43685;
  tmp_ivl_43693 <= fresh(293);
  LPM_q_ivl_43695 <= tmp_ivl_43697 & tmp_ivl_43693;
  new_AGEMA_signal_3268 <= tmp_ivl_43701(1);
  tmp_ivl_43699 <= tmp_ivl_43701(0);
  tmp_ivl_43701 <= LPM_d0_ivl_43705(0 + 1 downto 0);
  tmp_ivl_43706 <= new_AGEMA_signal_2963 & SboxInst_n323;
  LPM_q_ivl_43709 <= tmp_ivl_43711 & tmp_ivl_43706;
  tmp_ivl_43714 <= y4(7);
  tmp_ivl_43715 <= new_AGEMA_signal_2344 & tmp_ivl_43714;
  LPM_q_ivl_43718 <= tmp_ivl_43720 & tmp_ivl_43715;
  tmp_ivl_43723 <= fresh(294);
  LPM_q_ivl_43725 <= tmp_ivl_43727 & tmp_ivl_43723;
  new_AGEMA_signal_3269 <= tmp_ivl_43731(1);
  tmp_ivl_43729 <= tmp_ivl_43731(0);
  tmp_ivl_43731 <= LPM_d0_ivl_43735(0 + 1 downto 0);
  tmp_ivl_43736 <= new_AGEMA_signal_2964 & SboxInst_n376;
  LPM_q_ivl_43739 <= tmp_ivl_43741 & tmp_ivl_43736;
  tmp_ivl_43744 <= y4(17);
  tmp_ivl_43745 <= new_AGEMA_signal_2503 & tmp_ivl_43744;
  LPM_q_ivl_43748 <= tmp_ivl_43750 & tmp_ivl_43745;
  tmp_ivl_43753 <= fresh(295);
  LPM_q_ivl_43755 <= tmp_ivl_43757 & tmp_ivl_43753;
  new_AGEMA_signal_3270 <= tmp_ivl_43761(1);
  tmp_ivl_43759 <= tmp_ivl_43761(0);
  tmp_ivl_43761 <= LPM_d0_ivl_43765(0 + 1 downto 0);
  tmp_ivl_43766 <= new_AGEMA_signal_2965 & SboxInst_n368;
  LPM_q_ivl_43769 <= tmp_ivl_43771 & tmp_ivl_43766;
  tmp_ivl_43774 <= y4(24);
  tmp_ivl_43775 <= new_AGEMA_signal_2479 & tmp_ivl_43774;
  LPM_q_ivl_43778 <= tmp_ivl_43780 & tmp_ivl_43775;
  tmp_ivl_43783 <= fresh(296);
  LPM_q_ivl_43785 <= tmp_ivl_43787 & tmp_ivl_43783;
  new_AGEMA_signal_3271 <= tmp_ivl_43791(1);
  tmp_ivl_43789 <= tmp_ivl_43791(0);
  tmp_ivl_43791 <= LPM_d0_ivl_43795(0 + 1 downto 0);
  tmp_ivl_43796 <= new_AGEMA_signal_2966 & SboxInst_n324;
  LPM_q_ivl_43799 <= tmp_ivl_43801 & tmp_ivl_43796;
  tmp_ivl_43804 <= y4(6);
  tmp_ivl_43805 <= new_AGEMA_signal_2347 & tmp_ivl_43804;
  LPM_q_ivl_43808 <= tmp_ivl_43810 & tmp_ivl_43805;
  tmp_ivl_43813 <= fresh(297);
  LPM_q_ivl_43815 <= tmp_ivl_43817 & tmp_ivl_43813;
  new_AGEMA_signal_3272 <= tmp_ivl_43821(1);
  tmp_ivl_43819 <= tmp_ivl_43821(0);
  tmp_ivl_43821 <= LPM_d0_ivl_43825(0 + 1 downto 0);
  tmp_ivl_43826 <= new_AGEMA_signal_2967 & SboxInst_n369;
  LPM_q_ivl_43829 <= tmp_ivl_43831 & tmp_ivl_43826;
  tmp_ivl_43834 <= y4(23);
  tmp_ivl_43835 <= new_AGEMA_signal_2482 & tmp_ivl_43834;
  LPM_q_ivl_43838 <= tmp_ivl_43840 & tmp_ivl_43835;
  tmp_ivl_43843 <= fresh(298);
  LPM_q_ivl_43845 <= tmp_ivl_43847 & tmp_ivl_43843;
  new_AGEMA_signal_3273 <= tmp_ivl_43851(1);
  tmp_ivl_43849 <= tmp_ivl_43851(0);
  tmp_ivl_43851 <= LPM_d0_ivl_43855(0 + 1 downto 0);
  tmp_ivl_43856 <= new_AGEMA_signal_2968 & SboxInst_n377;
  LPM_q_ivl_43859 <= tmp_ivl_43861 & tmp_ivl_43856;
  tmp_ivl_43864 <= y4(16);
  tmp_ivl_43865 <= new_AGEMA_signal_2506 & tmp_ivl_43864;
  LPM_q_ivl_43868 <= tmp_ivl_43870 & tmp_ivl_43865;
  tmp_ivl_43873 <= fresh(299);
  LPM_q_ivl_43875 <= tmp_ivl_43877 & tmp_ivl_43873;
  new_AGEMA_signal_3274 <= tmp_ivl_43881(1);
  tmp_ivl_43879 <= tmp_ivl_43881(0);
  tmp_ivl_43881 <= LPM_d0_ivl_43885(0 + 1 downto 0);
  tmp_ivl_43886 <= new_AGEMA_signal_2969 & SboxInst_n370;
  LPM_q_ivl_43889 <= tmp_ivl_43891 & tmp_ivl_43886;
  tmp_ivl_43894 <= y4(22);
  tmp_ivl_43895 <= new_AGEMA_signal_2485 & tmp_ivl_43894;
  LPM_q_ivl_43898 <= tmp_ivl_43900 & tmp_ivl_43895;
  tmp_ivl_43903 <= fresh(300);
  LPM_q_ivl_43905 <= tmp_ivl_43907 & tmp_ivl_43903;
  new_AGEMA_signal_3275 <= tmp_ivl_43911(1);
  tmp_ivl_43909 <= tmp_ivl_43911(0);
  tmp_ivl_43911 <= LPM_d0_ivl_43915(0 + 1 downto 0);
  tmp_ivl_43916 <= new_AGEMA_signal_2970 & SboxInst_n378;
  LPM_q_ivl_43919 <= tmp_ivl_43921 & tmp_ivl_43916;
  tmp_ivl_43924 <= y4(15);
  tmp_ivl_43925 <= new_AGEMA_signal_2509 & tmp_ivl_43924;
  LPM_q_ivl_43928 <= tmp_ivl_43930 & tmp_ivl_43925;
  tmp_ivl_43933 <= fresh(301);
  LPM_q_ivl_43935 <= tmp_ivl_43937 & tmp_ivl_43933;
  new_AGEMA_signal_3276 <= tmp_ivl_43941(1);
  tmp_ivl_43939 <= tmp_ivl_43941(0);
  tmp_ivl_43941 <= LPM_d0_ivl_43945(0 + 1 downto 0);
  tmp_ivl_43946 <= new_AGEMA_signal_2971 & SboxInst_n379;
  LPM_q_ivl_43949 <= tmp_ivl_43951 & tmp_ivl_43946;
  tmp_ivl_43954 <= y4(14);
  tmp_ivl_43955 <= new_AGEMA_signal_2512 & tmp_ivl_43954;
  LPM_q_ivl_43958 <= tmp_ivl_43960 & tmp_ivl_43955;
  tmp_ivl_43963 <= fresh(302);
  LPM_q_ivl_43965 <= tmp_ivl_43967 & tmp_ivl_43963;
  new_AGEMA_signal_3277 <= tmp_ivl_43971(1);
  tmp_ivl_43969 <= tmp_ivl_43971(0);
  tmp_ivl_43971 <= LPM_d0_ivl_43975(0 + 1 downto 0);
  tmp_ivl_43976 <= new_AGEMA_signal_2972 & SboxInst_n371;
  LPM_q_ivl_43979 <= tmp_ivl_43981 & tmp_ivl_43976;
  tmp_ivl_43984 <= y4(21);
  tmp_ivl_43985 <= new_AGEMA_signal_2488 & tmp_ivl_43984;
  LPM_q_ivl_43988 <= tmp_ivl_43990 & tmp_ivl_43985;
  tmp_ivl_43993 <= fresh(303);
  LPM_q_ivl_43995 <= tmp_ivl_43997 & tmp_ivl_43993;
  new_AGEMA_signal_3278 <= tmp_ivl_44001(1);
  tmp_ivl_43999 <= tmp_ivl_44001(0);
  tmp_ivl_44001 <= LPM_d0_ivl_44005(0 + 1 downto 0);
  tmp_ivl_44006 <= new_AGEMA_signal_2973 & SboxInst_n372;
  LPM_q_ivl_44009 <= tmp_ivl_44011 & tmp_ivl_44006;
  tmp_ivl_44014 <= y4(20);
  tmp_ivl_44015 <= new_AGEMA_signal_2491 & tmp_ivl_44014;
  LPM_q_ivl_44018 <= tmp_ivl_44020 & tmp_ivl_44015;
  tmp_ivl_44023 <= fresh(304);
  LPM_q_ivl_44025 <= tmp_ivl_44027 & tmp_ivl_44023;
  new_AGEMA_signal_3279 <= tmp_ivl_44031(1);
  tmp_ivl_44029 <= tmp_ivl_44031(0);
  tmp_ivl_44031 <= LPM_d0_ivl_44035(0 + 1 downto 0);
  tmp_ivl_44036 <= new_AGEMA_signal_2974 & SboxInst_n380;
  LPM_q_ivl_44039 <= tmp_ivl_44041 & tmp_ivl_44036;
  tmp_ivl_44044 <= y4(13);
  tmp_ivl_44045 <= new_AGEMA_signal_2515 & tmp_ivl_44044;
  LPM_q_ivl_44048 <= tmp_ivl_44050 & tmp_ivl_44045;
  tmp_ivl_44053 <= fresh(305);
  LPM_q_ivl_44055 <= tmp_ivl_44057 & tmp_ivl_44053;
  new_AGEMA_signal_3280 <= tmp_ivl_44061(1);
  tmp_ivl_44059 <= tmp_ivl_44061(0);
  tmp_ivl_44061 <= LPM_d0_ivl_44065(0 + 1 downto 0);
  tmp_ivl_44066 <= new_AGEMA_signal_2975 & SboxInst_n381;
  LPM_q_ivl_44069 <= tmp_ivl_44071 & tmp_ivl_44066;
  tmp_ivl_44074 <= y4(12);
  tmp_ivl_44075 <= new_AGEMA_signal_2518 & tmp_ivl_44074;
  LPM_q_ivl_44078 <= tmp_ivl_44080 & tmp_ivl_44075;
  tmp_ivl_44083 <= fresh(306);
  LPM_q_ivl_44085 <= tmp_ivl_44087 & tmp_ivl_44083;
  new_AGEMA_signal_3281 <= tmp_ivl_44091(1);
  tmp_ivl_44089 <= tmp_ivl_44091(0);
  tmp_ivl_44091 <= LPM_d0_ivl_44095(0 + 1 downto 0);
  tmp_ivl_44096 <= new_AGEMA_signal_2976 & SboxInst_n374;
  LPM_q_ivl_44099 <= tmp_ivl_44101 & tmp_ivl_44096;
  tmp_ivl_44104 <= y4(19);
  tmp_ivl_44105 <= new_AGEMA_signal_2497 & tmp_ivl_44104;
  LPM_q_ivl_44108 <= tmp_ivl_44110 & tmp_ivl_44105;
  tmp_ivl_44113 <= fresh(307);
  LPM_q_ivl_44115 <= tmp_ivl_44117 & tmp_ivl_44113;
  new_AGEMA_signal_3282 <= tmp_ivl_44121(1);
  tmp_ivl_44119 <= tmp_ivl_44121(0);
  tmp_ivl_44121 <= LPM_d0_ivl_44125(0 + 1 downto 0);
  tmp_ivl_44126 <= new_AGEMA_signal_2977 & SboxInst_n382;
  LPM_q_ivl_44129 <= tmp_ivl_44131 & tmp_ivl_44126;
  tmp_ivl_44134 <= y4(11);
  tmp_ivl_44135 <= new_AGEMA_signal_2521 & tmp_ivl_44134;
  LPM_q_ivl_44138 <= tmp_ivl_44140 & tmp_ivl_44135;
  tmp_ivl_44143 <= fresh(308);
  LPM_q_ivl_44145 <= tmp_ivl_44147 & tmp_ivl_44143;
  new_AGEMA_signal_3283 <= tmp_ivl_44151(1);
  tmp_ivl_44149 <= tmp_ivl_44151(0);
  tmp_ivl_44151 <= LPM_d0_ivl_44155(0 + 1 downto 0);
  tmp_ivl_44156 <= new_AGEMA_signal_2978 & SboxInst_n375;
  LPM_q_ivl_44159 <= tmp_ivl_44161 & tmp_ivl_44156;
  tmp_ivl_44164 <= y4(18);
  tmp_ivl_44165 <= new_AGEMA_signal_2500 & tmp_ivl_44164;
  LPM_q_ivl_44168 <= tmp_ivl_44170 & tmp_ivl_44165;
  tmp_ivl_44173 <= fresh(309);
  LPM_q_ivl_44175 <= tmp_ivl_44177 & tmp_ivl_44173;
  new_AGEMA_signal_3284 <= tmp_ivl_44181(1);
  tmp_ivl_44179 <= tmp_ivl_44181(0);
  tmp_ivl_44181 <= LPM_d0_ivl_44185(0 + 1 downto 0);
  tmp_ivl_44186 <= new_AGEMA_signal_2979 & SboxInst_n383;
  LPM_q_ivl_44189 <= tmp_ivl_44191 & tmp_ivl_44186;
  tmp_ivl_44194 <= y4(10);
  tmp_ivl_44195 <= new_AGEMA_signal_2524 & tmp_ivl_44194;
  LPM_q_ivl_44198 <= tmp_ivl_44200 & tmp_ivl_44195;
  tmp_ivl_44203 <= fresh(310);
  LPM_q_ivl_44205 <= tmp_ivl_44207 & tmp_ivl_44203;
  new_AGEMA_signal_3285 <= tmp_ivl_44211(1);
  tmp_ivl_44209 <= tmp_ivl_44211(0);
  tmp_ivl_44211 <= LPM_d0_ivl_44215(0 + 1 downto 0);
  tmp_ivl_44216 <= new_AGEMA_signal_2980 & SboxInst_n367;
  LPM_q_ivl_44219 <= tmp_ivl_44221 & tmp_ivl_44216;
  tmp_ivl_44224 <= y4(25);
  tmp_ivl_44225 <= new_AGEMA_signal_2476 & tmp_ivl_44224;
  LPM_q_ivl_44228 <= tmp_ivl_44230 & tmp_ivl_44225;
  tmp_ivl_44233 <= fresh(311);
  LPM_q_ivl_44235 <= tmp_ivl_44237 & tmp_ivl_44233;
  new_AGEMA_signal_3286 <= tmp_ivl_44241(1);
  tmp_ivl_44239 <= tmp_ivl_44241(0);
  tmp_ivl_44241 <= LPM_d0_ivl_44245(0 + 1 downto 0);
  tmp_ivl_44246 <= new_AGEMA_signal_2981 & SboxInst_n360;
  LPM_q_ivl_44249 <= tmp_ivl_44251 & tmp_ivl_44246;
  tmp_ivl_44254 <= y4(31);
  tmp_ivl_44255 <= new_AGEMA_signal_2455 & tmp_ivl_44254;
  LPM_q_ivl_44258 <= tmp_ivl_44260 & tmp_ivl_44255;
  tmp_ivl_44263 <= fresh(312);
  LPM_q_ivl_44265 <= tmp_ivl_44267 & tmp_ivl_44263;
  new_AGEMA_signal_3287 <= tmp_ivl_44271(1);
  tmp_ivl_44269 <= tmp_ivl_44271(0);
  tmp_ivl_44271 <= LPM_d0_ivl_44275(0 + 1 downto 0);
  tmp_ivl_44276 <= new_AGEMA_signal_2982 & SboxInst_n361;
  LPM_q_ivl_44279 <= tmp_ivl_44281 & tmp_ivl_44276;
  tmp_ivl_44284 <= y4(30);
  tmp_ivl_44285 <= new_AGEMA_signal_2458 & tmp_ivl_44284;
  LPM_q_ivl_44288 <= tmp_ivl_44290 & tmp_ivl_44285;
  tmp_ivl_44293 <= fresh(313);
  LPM_q_ivl_44295 <= tmp_ivl_44297 & tmp_ivl_44293;
  new_AGEMA_signal_3288 <= tmp_ivl_44301(1);
  tmp_ivl_44299 <= tmp_ivl_44301(0);
  tmp_ivl_44301 <= LPM_d0_ivl_44305(0 + 1 downto 0);
  tmp_ivl_44306 <= new_AGEMA_signal_2983 & SboxInst_n363;
  LPM_q_ivl_44309 <= tmp_ivl_44311 & tmp_ivl_44306;
  tmp_ivl_44314 <= y4(29);
  tmp_ivl_44315 <= new_AGEMA_signal_2464 & tmp_ivl_44314;
  LPM_q_ivl_44318 <= tmp_ivl_44320 & tmp_ivl_44315;
  tmp_ivl_44323 <= fresh(314);
  LPM_q_ivl_44325 <= tmp_ivl_44327 & tmp_ivl_44323;
  new_AGEMA_signal_3289 <= tmp_ivl_44331(1);
  tmp_ivl_44329 <= tmp_ivl_44331(0);
  tmp_ivl_44331 <= LPM_d0_ivl_44335(0 + 1 downto 0);
  tmp_ivl_44336 <= new_AGEMA_signal_2984 & SboxInst_n364;
  LPM_q_ivl_44339 <= tmp_ivl_44341 & tmp_ivl_44336;
  tmp_ivl_44344 <= y4(28);
  tmp_ivl_44345 <= new_AGEMA_signal_2467 & tmp_ivl_44344;
  LPM_q_ivl_44348 <= tmp_ivl_44350 & tmp_ivl_44345;
  tmp_ivl_44353 <= fresh(315);
  LPM_q_ivl_44355 <= tmp_ivl_44357 & tmp_ivl_44353;
  new_AGEMA_signal_3290 <= tmp_ivl_44361(1);
  tmp_ivl_44359 <= tmp_ivl_44361(0);
  tmp_ivl_44361 <= LPM_d0_ivl_44365(0 + 1 downto 0);
  tmp_ivl_44366 <= new_AGEMA_signal_2985 & SboxInst_n365;
  LPM_q_ivl_44369 <= tmp_ivl_44371 & tmp_ivl_44366;
  tmp_ivl_44374 <= y4(27);
  tmp_ivl_44375 <= new_AGEMA_signal_2470 & tmp_ivl_44374;
  LPM_q_ivl_44378 <= tmp_ivl_44380 & tmp_ivl_44375;
  tmp_ivl_44383 <= fresh(316);
  LPM_q_ivl_44385 <= tmp_ivl_44387 & tmp_ivl_44383;
  new_AGEMA_signal_3291 <= tmp_ivl_44391(1);
  tmp_ivl_44389 <= tmp_ivl_44391(0);
  tmp_ivl_44391 <= LPM_d0_ivl_44395(0 + 1 downto 0);
  tmp_ivl_44396 <= new_AGEMA_signal_2986 & SboxInst_n321;
  LPM_q_ivl_44399 <= tmp_ivl_44401 & tmp_ivl_44396;
  tmp_ivl_44404 <= y4(9);
  tmp_ivl_44405 <= new_AGEMA_signal_2338 & tmp_ivl_44404;
  LPM_q_ivl_44408 <= tmp_ivl_44410 & tmp_ivl_44405;
  tmp_ivl_44413 <= fresh(317);
  LPM_q_ivl_44415 <= tmp_ivl_44417 & tmp_ivl_44413;
  new_AGEMA_signal_3292 <= tmp_ivl_44421(1);
  tmp_ivl_44419 <= tmp_ivl_44421(0);
  tmp_ivl_44421 <= LPM_d0_ivl_44425(0 + 1 downto 0);
  tmp_ivl_44426 <= new_AGEMA_signal_2987 & SboxInst_n366;
  LPM_q_ivl_44429 <= tmp_ivl_44431 & tmp_ivl_44426;
  tmp_ivl_44434 <= y4(26);
  tmp_ivl_44435 <= new_AGEMA_signal_2473 & tmp_ivl_44434;
  LPM_q_ivl_44438 <= tmp_ivl_44440 & tmp_ivl_44435;
  tmp_ivl_44443 <= fresh(318);
  LPM_q_ivl_44445 <= tmp_ivl_44447 & tmp_ivl_44443;
  new_AGEMA_signal_3293 <= tmp_ivl_44451(1);
  tmp_ivl_44449 <= tmp_ivl_44451(0);
  tmp_ivl_44451 <= LPM_d0_ivl_44455(0 + 1 downto 0);
  tmp_ivl_44456 <= new_AGEMA_signal_2988 & SboxInst_n322;
  LPM_q_ivl_44459 <= tmp_ivl_44461 & tmp_ivl_44456;
  tmp_ivl_44464 <= y4(8);
  tmp_ivl_44465 <= new_AGEMA_signal_2341 & tmp_ivl_44464;
  LPM_q_ivl_44468 <= tmp_ivl_44470 & tmp_ivl_44465;
  tmp_ivl_44473 <= fresh(319);
  LPM_q_ivl_44475 <= tmp_ivl_44477 & tmp_ivl_44473;
  new_AGEMA_signal_3294 <= tmp_ivl_44481(1);
  tmp_ivl_44479 <= tmp_ivl_44481(0);
  tmp_ivl_44481 <= LPM_d0_ivl_44485(0 + 1 downto 0);
  y4 <= tmp_ivl_138 & tmp_ivl_167 & tmp_ivl_196 & tmp_ivl_225 & tmp_ivl_283 & tmp_ivl_312 & tmp_ivl_341 & tmp_ivl_370 & tmp_ivl_399 & tmp_ivl_428 & tmp_ivl_457 & tmp_ivl_486 & tmp_ivl_515 & tmp_ivl_544 & tmp_ivl_602 & tmp_ivl_631 & tmp_ivl_660 & tmp_ivl_689 & tmp_ivl_718 & tmp_ivl_747 & tmp_ivl_776 & tmp_ivl_805 & tmp_ivl_834 & tmp_ivl_863 & tmp_ivl_921 & tmp_ivl_950 & tmp_ivl_979 & tmp_ivl_1008 & tmp_ivl_1037 & tmp_ivl_1066 & tmp_ivl_1095 & tmp_ivl_1124 & tmp_ivl_1153 & tmp_ivl_1182 & tmp_ivl_1240 & tmp_ivl_1269 & tmp_ivl_1298 & tmp_ivl_1327 & tmp_ivl_1356 & tmp_ivl_1385 & tmp_ivl_1414 & tmp_ivl_1443 & tmp_ivl_1472 & tmp_ivl_1501 & tmp_ivl_1559 & tmp_ivl_1588 & tmp_ivl_1617 & tmp_ivl_1646 & tmp_ivl_1675 & tmp_ivl_1704 & tmp_ivl_1733 & tmp_ivl_1762 & tmp_ivl_1791 & tmp_ivl_1820 & tmp_ivl_22 & tmp_ivl_51 & tmp_ivl_80 & tmp_ivl_109 & tmp_ivl_254 & tmp_ivl_573 & tmp_ivl_892 & tmp_ivl_1211 & tmp_ivl_1530 & tmp_ivl_1849;
  y0 <= tmp_ivl_1994 & tmp_ivl_2023 & tmp_ivl_2052 & tmp_ivl_2081 & tmp_ivl_2139 & tmp_ivl_2168 & tmp_ivl_2197 & tmp_ivl_2226 & tmp_ivl_2255 & tmp_ivl_2284 & tmp_ivl_2313 & tmp_ivl_2342 & tmp_ivl_2371 & tmp_ivl_2400 & tmp_ivl_2458 & tmp_ivl_2487 & tmp_ivl_2516 & tmp_ivl_2545 & tmp_ivl_2574 & tmp_ivl_2603 & tmp_ivl_2632 & tmp_ivl_2661 & tmp_ivl_2690 & tmp_ivl_2719 & tmp_ivl_2777 & tmp_ivl_2806 & tmp_ivl_2835 & tmp_ivl_2864 & tmp_ivl_2893 & tmp_ivl_2922 & tmp_ivl_2951 & tmp_ivl_2980 & tmp_ivl_3009 & tmp_ivl_3038 & tmp_ivl_3096 & tmp_ivl_3125 & tmp_ivl_3154 & tmp_ivl_3183 & tmp_ivl_3212 & tmp_ivl_3241 & tmp_ivl_3270 & tmp_ivl_3299 & tmp_ivl_3328 & tmp_ivl_3357 & tmp_ivl_3415 & tmp_ivl_3444 & tmp_ivl_3473 & tmp_ivl_3502 & tmp_ivl_3531 & tmp_ivl_3560 & tmp_ivl_3589 & tmp_ivl_3618 & tmp_ivl_3647 & tmp_ivl_3676 & tmp_ivl_1878 & tmp_ivl_1907 & tmp_ivl_1936 & tmp_ivl_1965 & tmp_ivl_2110 & tmp_ivl_2429 & tmp_ivl_2748 & tmp_ivl_3067 & tmp_ivl_3386 & tmp_ivl_3705;
  y2 <= tmp_ivl_5832 & tmp_ivl_5620;
  state_out_s1 <= tmp_ivl_13267 & tmp_ivl_9254 & tmp_ivl_8930 & tmp_ivl_8606 & tmp_ivl_8420 & tmp_ivl_8234 & tmp_ivl_8048 & tmp_ivl_13225 & tmp_ivl_7862 & tmp_ivl_10124 & tmp_ivl_9116 & tmp_ivl_8792 & tmp_ivl_25457 & tmp_ivl_23940 & tmp_ivl_22068 & tmp_ivl_20666 & tmp_ivl_19915 & tmp_ivl_18381 & tmp_ivl_17087 & tmp_ivl_15640 & tmp_ivl_13889 & tmp_ivl_24496 & tmp_ivl_22964 & tmp_ivl_21176 & tmp_ivl_10886 & tmp_ivl_19873 & tmp_ivl_17777 & tmp_ivl_16313 & tmp_ivl_14801 & tmp_ivl_13135 & tmp_ivl_12490 & tmp_ivl_11872 & tmp_ivl_21134 & tmp_ivl_10796 & tmp_ivl_9986 & tmp_ivl_9848 & tmp_ivl_9758 & tmp_ivl_9668 & tmp_ivl_9530 & tmp_ivl_9392 & tmp_ivl_11830 & tmp_ivl_19279 & tmp_ivl_25415 & tmp_ivl_23898 & tmp_ivl_22026 & tmp_ivl_20624 & tmp_ivl_24454 & tmp_ivl_22922 & tmp_ivl_17045 & tmp_ivl_15598 & tmp_ivl_19831 & tmp_ivl_25373 & tmp_ivl_23856 & tmp_ivl_21984 & tmp_ivl_20582 & tmp_ivl_12448 & tmp_ivl_18339 & tmp_ivl_17003 & tmp_ivl_15556 & tmp_ivl_13847 & tmp_ivl_12580 & tmp_ivl_12161 & tmp_ivl_11024 & tmp_ivl_18297 & tmp_ivl_31816 & tmp_ivl_34531 & tmp_ivl_34701 & tmp_ivl_34913 & tmp_ivl_35041 & tmp_ivl_31457 & tmp_ivl_31266 & tmp_ivl_30479 & tmp_ivl_27116 & tmp_ivl_26879 & tmp_ivl_26642 & tmp_ivl_26405 & tmp_ivl_26168 & tmp_ivl_25931 & tmp_ivl_25694 & tmp_ivl_30586 & tmp_ivl_28167 & tmp_ivl_28060 & tmp_ivl_27953 & tmp_ivl_27846 & tmp_ivl_27739 & tmp_ivl_27632 & tmp_ivl_27460 & tmp_ivl_27288 & tmp_ivl_29023 & tmp_ivl_28916 & tmp_ivl_28809 & tmp_ivl_28702 & tmp_ivl_28595 & tmp_ivl_28488 & tmp_ivl_28381 & tmp_ivl_28274 & tmp_ivl_29879 & tmp_ivl_29772 & tmp_ivl_29665 & tmp_ivl_29558 & tmp_ivl_29451 & tmp_ivl_29344 & tmp_ivl_29237 & tmp_ivl_29130 & tmp_ivl_30437 & tmp_ivl_31054 & tmp_ivl_30842 & tmp_ivl_30693 & tmp_ivl_30307 & tmp_ivl_30200 & tmp_ivl_30093 & tmp_ivl_29986 & tmp_ivl_31224 & tmp_ivl_31774 & tmp_ivl_34573 & tmp_ivl_34743 & tmp_ivl_34871 & tmp_ivl_35083 & tmp_ivl_31415 & tmp_ivl_31182 & tmp_ivl_31012 & tmp_ivl_30800 & tmp_ivl_31732 & tmp_ivl_34615 & tmp_ivl_34785 & tmp_ivl_34955 & tmp_ivl_35125 & tmp_ivl_31373 & tmp_ivl_34109 & tmp_ivl_31646 & tmp_ivl_34172 & tmp_ivl_34235 & tmp_ivl_34277 & tmp_ivl_31562 & tmp_ivl_34361 & tmp_ivl_31967 & tmp_ivl_33773 & tmp_ivl_33815 & tmp_ivl_33857 & tmp_ivl_33899 & tmp_ivl_33941 & tmp_ivl_33983 & tmp_ivl_34025 & tmp_ivl_34067 & tmp_ivl_33437 & tmp_ivl_33479 & tmp_ivl_33521 & tmp_ivl_33563 & tmp_ivl_33605 & tmp_ivl_33647 & tmp_ivl_33689 & tmp_ivl_33731 & tmp_ivl_33101 & tmp_ivl_33143 & tmp_ivl_33185 & tmp_ivl_33227 & tmp_ivl_33269 & tmp_ivl_33311 & tmp_ivl_33353 & tmp_ivl_33395 & tmp_ivl_32765 & tmp_ivl_32807 & tmp_ivl_32849 & tmp_ivl_32891 & tmp_ivl_32933 & tmp_ivl_32975 & tmp_ivl_33017 & tmp_ivl_33059 & tmp_ivl_32429 & tmp_ivl_32471 & tmp_ivl_32513 & tmp_ivl_32555 & tmp_ivl_32597 & tmp_ivl_32639 & tmp_ivl_32681 & tmp_ivl_32723 & tmp_ivl_32093 & tmp_ivl_32135 & tmp_ivl_32177 & tmp_ivl_32219 & tmp_ivl_32261 & tmp_ivl_32303 & tmp_ivl_32345 & tmp_ivl_32387 & tmp_ivl_31902 & tmp_ivl_30926 & tmp_ivl_31520 & tmp_ivl_34319 & tmp_ivl_34403 & tmp_ivl_34445 & tmp_ivl_32009 & tmp_ivl_32051 & tmp_ivl_25138 & tmp_ivl_23621 & tmp_ivl_22431 & tmp_ivl_25096 & tmp_ivl_23579 & tmp_ivl_21791 & tmp_ivl_20945 & tmp_ivl_20194 & tmp_ivl_17370 & tmp_ivl_16057 & tmp_ivl_15151 & tmp_ivl_16913 & tmp_ivl_15466 & tmp_ivl_24775 & tmp_ivl_22710 & tmp_ivl_22389 & tmp_ivl_18748 & tmp_ivl_17993 & tmp_ivl_11514 & tmp_ivl_12071 & tmp_ivl_11740 & tmp_ivl_16571 & tmp_ivl_15774 & tmp_ivl_14562 & tmp_ivl_22668 & tmp_ivl_22347 & tmp_ivl_25054 & tmp_ivl_23537 & tmp_ivl_21749 & tmp_ivl_20903 & tmp_ivl_20152 & tmp_ivl_19090 & tmp_ivl_17584 & tmp_ivl_14520 & tmp_ivl_16871 & tmp_ivl_15424 & tmp_ivl_14195 & tmp_ivl_13493 & tmp_ivl_12806 & tmp_ivl_24733 & tmp_ivl_21470 & tmp_ivl_24219 & tmp_ivl_23258 & tmp_ivl_21428 & tmp_ivl_20389 & tmp_ivl_19680 & tmp_ivl_19466 & tmp_ivl_18207 & tmp_ivl_15109 & tmp_ivl_17328 & tmp_ivl_16015 & tmp_ivl_15067 & tmp_ivl_13757 & tmp_ivl_13045 & tmp_ivl_24177 & tmp_ivl_23216 & tmp_ivl_18981 & tmp_ivl_18614 & tmp_ivl_17911 & tmp_ivl_11315 & tmp_ivl_10706 & tmp_ivl_10415 & tmp_ivl_17221 & tmp_ivl_15908 & tmp_ivl_24624 & tmp_ivl_22559 & tmp_ivl_22238 & tmp_ivl_24945 & tmp_ivl_23428 & tmp_ivl_21640 & tmp_ivl_20794 & tmp_ivl_20043 & tmp_ivl_20280 & tmp_ivl_19571 & tmp_ivl_19384 & tmp_ivl_18098 & tmp_ivl_19766 & tmp_ivl_17712 & tmp_ivl_16248 & tmp_ivl_14736 & tmp_ivl_23791 & tmp_ivl_21919 & tmp_ivl_20517 & tmp_ivl_17475 & tmp_ivl_12310 & tmp_ivl_24389 & tmp_ivl_23134 & tmp_ivl_21346 & tmp_ivl_21877 & tmp_ivl_20475 & tmp_ivl_17670 & tmp_ivl_16143 & tmp_ivl_24068 & tmp_ivl_23092 & tmp_ivl_21304 & tmp_ivl_25308 & tmp_ivl_23386 & tmp_ivl_21598 & tmp_ivl_20752 & tmp_ivl_20001 & tmp_ivl_18872 & tmp_ivl_18505 & tmp_ivl_25266 & tmp_ivl_23749 & tmp_ivl_21556 & tmp_ivl_24026 & tmp_ivl_23050 & tmp_ivl_21262 & tmp_ivl_24582 & tmp_ivl_22517 & tmp_ivl_22196 & tmp_ivl_24903 & tmp_ivl_13994 & tmp_ivl_24347 & tmp_ivl_22857 & tmp_ivl_25224 & tmp_ivl_23707 & tmp_ivl_22154 & tmp_ivl_24861 & tmp_ivl_23344 & tmp_ivl_24305 & tmp_ivl_22815 & tmp_ivl_21069 & tmp_ivl_16462 & tmp_ivl_19214 & tmp_ivl_14344 & tmp_ivl_16695 & tmp_ivl_15275;
  state_out_s0 <= tmp_ivl_13269 & tmp_ivl_9256 & tmp_ivl_8932 & tmp_ivl_8608 & tmp_ivl_8422 & tmp_ivl_8236 & tmp_ivl_8050 & tmp_ivl_13227 & tmp_ivl_7864 & tmp_ivl_10126 & tmp_ivl_9118 & tmp_ivl_8794 & tmp_ivl_25459 & tmp_ivl_23942 & tmp_ivl_22070 & tmp_ivl_20668 & tmp_ivl_19917 & tmp_ivl_18383 & tmp_ivl_17089 & tmp_ivl_15642 & tmp_ivl_13891 & tmp_ivl_24498 & tmp_ivl_22966 & tmp_ivl_21178 & tmp_ivl_10888 & tmp_ivl_19875 & tmp_ivl_17779 & tmp_ivl_16315 & tmp_ivl_14803 & tmp_ivl_13137 & tmp_ivl_12492 & tmp_ivl_11874 & tmp_ivl_21136 & tmp_ivl_10798 & tmp_ivl_9988 & tmp_ivl_9850 & tmp_ivl_9760 & tmp_ivl_9670 & tmp_ivl_9532 & tmp_ivl_9394 & tmp_ivl_11832 & tmp_ivl_19281 & tmp_ivl_25417 & tmp_ivl_23900 & tmp_ivl_22028 & tmp_ivl_20626 & tmp_ivl_24456 & tmp_ivl_22924 & tmp_ivl_17047 & tmp_ivl_15600 & tmp_ivl_19833 & tmp_ivl_25375 & tmp_ivl_23858 & tmp_ivl_21986 & tmp_ivl_20584 & tmp_ivl_12450 & tmp_ivl_18341 & tmp_ivl_17005 & tmp_ivl_15558 & tmp_ivl_13849 & tmp_ivl_12582 & tmp_ivl_12163 & tmp_ivl_11026 & tmp_ivl_18299 & tmp_ivl_31818 & tmp_ivl_34533 & tmp_ivl_34703 & tmp_ivl_34915 & tmp_ivl_35043 & tmp_ivl_31459 & tmp_ivl_31268 & tmp_ivl_30481 & tmp_ivl_27118 & tmp_ivl_26881 & tmp_ivl_26644 & tmp_ivl_26407 & tmp_ivl_26170 & tmp_ivl_25933 & tmp_ivl_25696 & tmp_ivl_30588 & tmp_ivl_28169 & tmp_ivl_28062 & tmp_ivl_27955 & tmp_ivl_27848 & tmp_ivl_27741 & tmp_ivl_27634 & tmp_ivl_27462 & tmp_ivl_27290 & tmp_ivl_29025 & tmp_ivl_28918 & tmp_ivl_28811 & tmp_ivl_28704 & tmp_ivl_28597 & tmp_ivl_28490 & tmp_ivl_28383 & tmp_ivl_28276 & tmp_ivl_29881 & tmp_ivl_29774 & tmp_ivl_29667 & tmp_ivl_29560 & tmp_ivl_29453 & tmp_ivl_29346 & tmp_ivl_29239 & tmp_ivl_29132 & tmp_ivl_30439 & tmp_ivl_31056 & tmp_ivl_30844 & tmp_ivl_30695 & tmp_ivl_30309 & tmp_ivl_30202 & tmp_ivl_30095 & tmp_ivl_29988 & tmp_ivl_31226 & tmp_ivl_31776 & tmp_ivl_34575 & tmp_ivl_34745 & tmp_ivl_34873 & tmp_ivl_35085 & tmp_ivl_31417 & tmp_ivl_31184 & tmp_ivl_31014 & tmp_ivl_30802 & tmp_ivl_31734 & tmp_ivl_34617 & tmp_ivl_34787 & tmp_ivl_34957 & tmp_ivl_35127 & tmp_ivl_31375 & tmp_ivl_34111 & tmp_ivl_31648 & tmp_ivl_34174 & tmp_ivl_34237 & tmp_ivl_34279 & tmp_ivl_31564 & tmp_ivl_34363 & tmp_ivl_31969 & tmp_ivl_33775 & tmp_ivl_33817 & tmp_ivl_33859 & tmp_ivl_33901 & tmp_ivl_33943 & tmp_ivl_33985 & tmp_ivl_34027 & tmp_ivl_34069 & tmp_ivl_33439 & tmp_ivl_33481 & tmp_ivl_33523 & tmp_ivl_33565 & tmp_ivl_33607 & tmp_ivl_33649 & tmp_ivl_33691 & tmp_ivl_33733 & tmp_ivl_33103 & tmp_ivl_33145 & tmp_ivl_33187 & tmp_ivl_33229 & tmp_ivl_33271 & tmp_ivl_33313 & tmp_ivl_33355 & tmp_ivl_33397 & tmp_ivl_32767 & tmp_ivl_32809 & tmp_ivl_32851 & tmp_ivl_32893 & tmp_ivl_32935 & tmp_ivl_32977 & tmp_ivl_33019 & tmp_ivl_33061 & tmp_ivl_32431 & tmp_ivl_32473 & tmp_ivl_32515 & tmp_ivl_32557 & tmp_ivl_32599 & tmp_ivl_32641 & tmp_ivl_32683 & tmp_ivl_32725 & tmp_ivl_32095 & tmp_ivl_32137 & tmp_ivl_32179 & tmp_ivl_32221 & tmp_ivl_32263 & tmp_ivl_32305 & tmp_ivl_32347 & tmp_ivl_32389 & tmp_ivl_31904 & tmp_ivl_30928 & tmp_ivl_31522 & tmp_ivl_34321 & tmp_ivl_34405 & tmp_ivl_34447 & tmp_ivl_32011 & tmp_ivl_32053 & tmp_ivl_25140 & tmp_ivl_23623 & tmp_ivl_22433 & tmp_ivl_25098 & tmp_ivl_23581 & tmp_ivl_21793 & tmp_ivl_20947 & tmp_ivl_20196 & tmp_ivl_17372 & tmp_ivl_16059 & tmp_ivl_15153 & tmp_ivl_16915 & tmp_ivl_15468 & tmp_ivl_24777 & tmp_ivl_22712 & tmp_ivl_22391 & tmp_ivl_18750 & tmp_ivl_17995 & tmp_ivl_11516 & tmp_ivl_12073 & tmp_ivl_11742 & tmp_ivl_16573 & tmp_ivl_15776 & tmp_ivl_14564 & tmp_ivl_22670 & tmp_ivl_22349 & tmp_ivl_25056 & tmp_ivl_23539 & tmp_ivl_21751 & tmp_ivl_20905 & tmp_ivl_20154 & tmp_ivl_19092 & tmp_ivl_17586 & tmp_ivl_14522 & tmp_ivl_16873 & tmp_ivl_15426 & tmp_ivl_14197 & tmp_ivl_13495 & tmp_ivl_12808 & tmp_ivl_24735 & tmp_ivl_21472 & tmp_ivl_24221 & tmp_ivl_23260 & tmp_ivl_21430 & tmp_ivl_20391 & tmp_ivl_19682 & tmp_ivl_19468 & tmp_ivl_18209 & tmp_ivl_15111 & tmp_ivl_17330 & tmp_ivl_16017 & tmp_ivl_15069 & tmp_ivl_13759 & tmp_ivl_13047 & tmp_ivl_24179 & tmp_ivl_23218 & tmp_ivl_18983 & tmp_ivl_18616 & tmp_ivl_17913 & tmp_ivl_11317 & tmp_ivl_10708 & tmp_ivl_10417 & tmp_ivl_17223 & tmp_ivl_15910 & tmp_ivl_24626 & tmp_ivl_22561 & tmp_ivl_22240 & tmp_ivl_24947 & tmp_ivl_23430 & tmp_ivl_21642 & tmp_ivl_20796 & tmp_ivl_20045 & tmp_ivl_20282 & tmp_ivl_19573 & tmp_ivl_19386 & tmp_ivl_18100 & tmp_ivl_19768 & tmp_ivl_17714 & tmp_ivl_16250 & tmp_ivl_14738 & tmp_ivl_23793 & tmp_ivl_21921 & tmp_ivl_20519 & tmp_ivl_17477 & tmp_ivl_12312 & tmp_ivl_24391 & tmp_ivl_23136 & tmp_ivl_21348 & tmp_ivl_21879 & tmp_ivl_20477 & tmp_ivl_17672 & tmp_ivl_16145 & tmp_ivl_24070 & tmp_ivl_23094 & tmp_ivl_21306 & tmp_ivl_25310 & tmp_ivl_23388 & tmp_ivl_21600 & tmp_ivl_20754 & tmp_ivl_20003 & tmp_ivl_18874 & tmp_ivl_18507 & tmp_ivl_25268 & tmp_ivl_23751 & tmp_ivl_21558 & tmp_ivl_24028 & tmp_ivl_23052 & tmp_ivl_21264 & tmp_ivl_24584 & tmp_ivl_22519 & tmp_ivl_22198 & tmp_ivl_24905 & tmp_ivl_13996 & tmp_ivl_24349 & tmp_ivl_22859 & tmp_ivl_25226 & tmp_ivl_23709 & tmp_ivl_22156 & tmp_ivl_24863 & tmp_ivl_23346 & tmp_ivl_24307 & tmp_ivl_22817 & tmp_ivl_21071 & tmp_ivl_16464 & tmp_ivl_19216 & tmp_ivl_14346 & tmp_ivl_16697 & tmp_ivl_15277;
  z1 <= tmp_ivl_36811 & tmp_ivl_36783 & tmp_ivl_36755 & tmp_ivl_36727 & tmp_ivl_36671 & tmp_ivl_36643 & tmp_ivl_36615 & tmp_ivl_36587 & tmp_ivl_36559 & tmp_ivl_36531 & tmp_ivl_36503 & tmp_ivl_36475 & tmp_ivl_36447 & tmp_ivl_36419 & tmp_ivl_36363 & tmp_ivl_36335 & tmp_ivl_36307 & tmp_ivl_36279 & tmp_ivl_36251 & tmp_ivl_36223 & tmp_ivl_36195 & tmp_ivl_36167 & tmp_ivl_36139 & tmp_ivl_36111 & tmp_ivl_36055 & tmp_ivl_36027 & tmp_ivl_35999 & tmp_ivl_35971 & tmp_ivl_35943 & tmp_ivl_35915 & tmp_ivl_35887 & tmp_ivl_35859 & tmp_ivl_35831 & tmp_ivl_35803 & tmp_ivl_35747 & tmp_ivl_35719 & tmp_ivl_35691 & tmp_ivl_35663 & tmp_ivl_35635 & tmp_ivl_35607 & tmp_ivl_35579 & tmp_ivl_35551 & tmp_ivl_35523 & tmp_ivl_35495 & tmp_ivl_35437 & tmp_ivl_35409 & tmp_ivl_35381 & tmp_ivl_35353 & tmp_ivl_35325 & tmp_ivl_35297 & tmp_ivl_35269 & tmp_ivl_35241 & tmp_ivl_35213 & tmp_ivl_35185 & tmp_ivl_36923 & tmp_ivl_36895 & tmp_ivl_36867 & tmp_ivl_36839 & tmp_ivl_36699 & tmp_ivl_36391 & tmp_ivl_36083 & tmp_ivl_35775 & tmp_ivl_35467 & tmp_ivl_35157;
  z3 <= tmp_ivl_38723 & tmp_ivl_38693 & tmp_ivl_38663 & tmp_ivl_38633 & tmp_ivl_38573 & tmp_ivl_38543 & tmp_ivl_38513 & tmp_ivl_38483 & tmp_ivl_38453 & tmp_ivl_38423 & tmp_ivl_38393 & tmp_ivl_38363 & tmp_ivl_38333 & tmp_ivl_38303 & tmp_ivl_38243 & tmp_ivl_38213 & tmp_ivl_38183 & tmp_ivl_38153 & tmp_ivl_38123 & tmp_ivl_38093 & tmp_ivl_38063 & tmp_ivl_38033 & tmp_ivl_38003 & tmp_ivl_37973 & tmp_ivl_37913 & tmp_ivl_37883 & tmp_ivl_37853 & tmp_ivl_37823 & tmp_ivl_37793 & tmp_ivl_37763 & tmp_ivl_37733 & tmp_ivl_37703 & tmp_ivl_37673 & tmp_ivl_37643 & tmp_ivl_37583 & tmp_ivl_37553 & tmp_ivl_37523 & tmp_ivl_37493 & tmp_ivl_37463 & tmp_ivl_37433 & tmp_ivl_37403 & tmp_ivl_37373 & tmp_ivl_37343 & tmp_ivl_37313 & tmp_ivl_37253 & tmp_ivl_37223 & tmp_ivl_37193 & tmp_ivl_37163 & tmp_ivl_37133 & tmp_ivl_37103 & tmp_ivl_37073 & tmp_ivl_37043 & tmp_ivl_37013 & tmp_ivl_36983 & tmp_ivl_38843 & tmp_ivl_38813 & tmp_ivl_38783 & tmp_ivl_38753 & tmp_ivl_38603 & tmp_ivl_38273 & tmp_ivl_37943 & tmp_ivl_37613 & tmp_ivl_37283 & tmp_ivl_36953;
  z4 <= tmp_ivl_40643 & tmp_ivl_40613 & tmp_ivl_40583 & tmp_ivl_40553 & tmp_ivl_40493 & tmp_ivl_40463 & tmp_ivl_40433 & tmp_ivl_40403 & tmp_ivl_40373 & tmp_ivl_40343 & tmp_ivl_40313 & tmp_ivl_40283 & tmp_ivl_40253 & tmp_ivl_40223 & tmp_ivl_40163 & tmp_ivl_40133 & tmp_ivl_40103 & tmp_ivl_40073 & tmp_ivl_40043 & tmp_ivl_40013 & tmp_ivl_39983 & tmp_ivl_39953 & tmp_ivl_39923 & tmp_ivl_39893 & tmp_ivl_39833 & tmp_ivl_39803 & tmp_ivl_39773 & tmp_ivl_39743 & tmp_ivl_39713 & tmp_ivl_39683 & tmp_ivl_39653 & tmp_ivl_39623 & tmp_ivl_39593 & tmp_ivl_39563 & tmp_ivl_39503 & tmp_ivl_39473 & tmp_ivl_39443 & tmp_ivl_39413 & tmp_ivl_39383 & tmp_ivl_39353 & tmp_ivl_39323 & tmp_ivl_39293 & tmp_ivl_39263 & tmp_ivl_39233 & tmp_ivl_39173 & tmp_ivl_39143 & tmp_ivl_39113 & tmp_ivl_39083 & tmp_ivl_39053 & tmp_ivl_39023 & tmp_ivl_38993 & tmp_ivl_38963 & tmp_ivl_38933 & tmp_ivl_38903 & tmp_ivl_40763 & tmp_ivl_40733 & tmp_ivl_40703 & tmp_ivl_40673 & tmp_ivl_40523 & tmp_ivl_40193 & tmp_ivl_39863 & tmp_ivl_39533 & tmp_ivl_39203 & tmp_ivl_38873;
  z2 <= tmp_ivl_41693 & tmp_ivl_41813 & tmp_ivl_41483 & tmp_ivl_41573 & tmp_ivl_41603 & tmp_ivl_41633 & tmp_ivl_41663 & tmp_ivl_41513 & tmp_ivl_41453 & tmp_ivl_41543 & tmp_ivl_41243 & tmp_ivl_41303 & tmp_ivl_41363 & tmp_ivl_41393 & tmp_ivl_41423 & tmp_ivl_41213 & tmp_ivl_41273 & tmp_ivl_41333 & tmp_ivl_40793 & tmp_ivl_40883 & tmp_ivl_40943 & tmp_ivl_41003 & tmp_ivl_41063 & tmp_ivl_40853 & tmp_ivl_40823 & tmp_ivl_40913 & tmp_ivl_40973 & tmp_ivl_41033 & tmp_ivl_41093 & tmp_ivl_41123 & tmp_ivl_41153 & tmp_ivl_41183 & tmp_ivl_44269 & tmp_ivl_44299 & tmp_ivl_44329 & tmp_ivl_44359 & tmp_ivl_44389 & tmp_ivl_44449 & tmp_ivl_44239 & tmp_ivl_43789 & tmp_ivl_43849 & tmp_ivl_43909 & tmp_ivl_43999 & tmp_ivl_44029 & tmp_ivl_44119 & tmp_ivl_44179 & tmp_ivl_43759 & tmp_ivl_43879 & tmp_ivl_43939 & tmp_ivl_43969 & tmp_ivl_44059 & tmp_ivl_44089 & tmp_ivl_44149 & tmp_ivl_44209 & tmp_ivl_44419 & tmp_ivl_44479 & tmp_ivl_43729 & tmp_ivl_43819 & tmp_ivl_41753 & tmp_ivl_41783 & tmp_ivl_41843 & tmp_ivl_41873 & tmp_ivl_41903 & tmp_ivl_41723;
  z0 <= tmp_ivl_42299 & tmp_ivl_42383 & tmp_ivl_42439 & tmp_ivl_43027 & tmp_ivl_43111 & tmp_ivl_43167 & tmp_ivl_43223 & tmp_ivl_43251 & tmp_ivl_43279 & tmp_ivl_42523 & tmp_ivl_42607 & tmp_ivl_42691 & tmp_ivl_42747 & tmp_ivl_42803 & tmp_ivl_42831 & tmp_ivl_42859 & tmp_ivl_42887 & tmp_ivl_41931 & tmp_ivl_42043 & tmp_ivl_42099 & tmp_ivl_42183 & tmp_ivl_42241 & tmp_ivl_42327 & tmp_ivl_42355 & tmp_ivl_42411 & tmp_ivl_43587 & tmp_ivl_43643 & tmp_ivl_43531 & tmp_ivl_43559 & tmp_ivl_43615 & tmp_ivl_43671 & tmp_ivl_43699 & tmp_ivl_43307 & tmp_ivl_43363 & tmp_ivl_43447 & tmp_ivl_43335 & tmp_ivl_43391 & tmp_ivl_43419 & tmp_ivl_43475 & tmp_ivl_43503 & tmp_ivl_42943 & tmp_ivl_42999 & tmp_ivl_43055 & tmp_ivl_42915 & tmp_ivl_42971 & tmp_ivl_43083 & tmp_ivl_43139 & tmp_ivl_43195 & tmp_ivl_42467 & tmp_ivl_42579 & tmp_ivl_42663 & tmp_ivl_42495 & tmp_ivl_42551 & tmp_ivl_42635 & tmp_ivl_42719 & tmp_ivl_42775 & tmp_ivl_41959 & tmp_ivl_42015 & tmp_ivl_42155 & tmp_ivl_41987 & tmp_ivl_42071 & tmp_ivl_42127 & tmp_ivl_42213 & tmp_ivl_42271;
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3355
  SboxInst_U1: not_masked
    port map (
      a => LPM_q_ivl_7681,
      b => LPM_d0_ivl_7683
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4945
  SboxInst_U10: and_HPC2
    port map (
      a => LPM_q_ivl_44339,
      b => LPM_q_ivl_44348,
      c => LPM_d0_ivl_44365,
      clk => clk,
      r => LPM_q_ivl_44355
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4900
  SboxInst_U100: and_HPC2
    port map (
      a => LPM_q_ivl_43037,
      b => LPM_q_ivl_43044,
      c => LPM_d0_ivl_43061,
      clk => clk,
      r => LPM_q_ivl_43051
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3305
  SboxInst_U101: not_masked
    port map (
      a => LPM_q_ivl_7231,
      b => LPM_d0_ivl_7233
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4899
  SboxInst_U102: and_HPC2
    port map (
      a => LPM_q_ivl_43009,
      b => LPM_q_ivl_43016,
      c => LPM_d0_ivl_43033,
      clk => clk,
      r => LPM_q_ivl_43023
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3304
  SboxInst_U103: not_masked
    port map (
      a => LPM_q_ivl_7222,
      b => LPM_d0_ivl_7224
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4898
  SboxInst_U104: and_HPC2
    port map (
      a => LPM_q_ivl_42981,
      b => LPM_q_ivl_42988,
      c => LPM_d0_ivl_43005,
      clk => clk,
      r => LPM_q_ivl_42995
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3303
  SboxInst_U105: not_masked
    port map (
      a => LPM_q_ivl_7213,
      b => LPM_d0_ivl_7215
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4897
  SboxInst_U106: and_HPC2
    port map (
      a => LPM_q_ivl_42953,
      b => LPM_q_ivl_42960,
      c => LPM_d0_ivl_42977,
      clk => clk,
      r => LPM_q_ivl_42967
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3302
  SboxInst_U107: not_masked
    port map (
      a => LPM_q_ivl_7204,
      b => LPM_d0_ivl_7206
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4896
  SboxInst_U108: and_HPC2
    port map (
      a => LPM_q_ivl_42925,
      b => LPM_q_ivl_42932,
      c => LPM_d0_ivl_42949,
      clk => clk,
      r => LPM_q_ivl_42939
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3301
  SboxInst_U109: not_masked
    port map (
      a => LPM_q_ivl_7195,
      b => LPM_d0_ivl_7197
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3350
  SboxInst_U11: not_masked
    port map (
      a => LPM_q_ivl_7636,
      b => LPM_d0_ivl_7638
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4895
  SboxInst_U110: and_HPC2
    port map (
      a => LPM_q_ivl_42897,
      b => LPM_q_ivl_42904,
      c => LPM_d0_ivl_42921,
      clk => clk,
      r => LPM_q_ivl_42911
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3300
  SboxInst_U111: not_masked
    port map (
      a => LPM_q_ivl_7186,
      b => LPM_d0_ivl_7188
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4894
  SboxInst_U112: and_HPC2
    port map (
      a => LPM_q_ivl_42869,
      b => LPM_q_ivl_42876,
      c => LPM_d0_ivl_42893,
      clk => clk,
      r => LPM_q_ivl_42883
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3299
  SboxInst_U113: not_masked
    port map (
      a => LPM_q_ivl_7177,
      b => LPM_d0_ivl_7179
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4893
  SboxInst_U114: and_HPC2
    port map (
      a => LPM_q_ivl_42841,
      b => LPM_q_ivl_42848,
      c => LPM_d0_ivl_42865,
      clk => clk,
      r => LPM_q_ivl_42855
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3298
  SboxInst_U115: not_masked
    port map (
      a => LPM_q_ivl_7168,
      b => LPM_d0_ivl_7170
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4892
  SboxInst_U116: and_HPC2
    port map (
      a => LPM_q_ivl_42813,
      b => LPM_q_ivl_42820,
      c => LPM_d0_ivl_42837,
      clk => clk,
      r => LPM_q_ivl_42827
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3297
  SboxInst_U117: not_masked
    port map (
      a => LPM_q_ivl_7159,
      b => LPM_d0_ivl_7161
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4891
  SboxInst_U118: and_HPC2
    port map (
      a => LPM_q_ivl_42785,
      b => LPM_q_ivl_42792,
      c => LPM_d0_ivl_42809,
      clk => clk,
      r => LPM_q_ivl_42799
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3296
  SboxInst_U119: not_masked
    port map (
      a => LPM_q_ivl_7150,
      b => LPM_d0_ivl_7152
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4944
  SboxInst_U12: and_HPC2
    port map (
      a => LPM_q_ivl_44309,
      b => LPM_q_ivl_44318,
      c => LPM_d0_ivl_44335,
      clk => clk,
      r => LPM_q_ivl_44325
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4890
  SboxInst_U120: and_HPC2
    port map (
      a => LPM_q_ivl_42757,
      b => LPM_q_ivl_42764,
      c => LPM_d0_ivl_42781,
      clk => clk,
      r => LPM_q_ivl_42771
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3295
  SboxInst_U121: not_masked
    port map (
      a => LPM_q_ivl_7141,
      b => LPM_d0_ivl_7143
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4889
  SboxInst_U122: and_HPC2
    port map (
      a => LPM_q_ivl_42729,
      b => LPM_q_ivl_42736,
      c => LPM_d0_ivl_42753,
      clk => clk,
      r => LPM_q_ivl_42743
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3294
  SboxInst_U123: not_masked
    port map (
      a => LPM_q_ivl_7132,
      b => LPM_d0_ivl_7134
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4888
  SboxInst_U124: and_HPC2
    port map (
      a => LPM_q_ivl_42701,
      b => LPM_q_ivl_42708,
      c => LPM_d0_ivl_42725,
      clk => clk,
      r => LPM_q_ivl_42715
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3293
  SboxInst_U125: not_masked
    port map (
      a => LPM_q_ivl_7123,
      b => LPM_d0_ivl_7125
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4887
  SboxInst_U126: and_HPC2
    port map (
      a => LPM_q_ivl_42673,
      b => LPM_q_ivl_42680,
      c => LPM_d0_ivl_42697,
      clk => clk,
      r => LPM_q_ivl_42687
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3292
  SboxInst_U127: not_masked
    port map (
      a => LPM_q_ivl_7114,
      b => LPM_d0_ivl_7116
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4886
  SboxInst_U128: and_HPC2
    port map (
      a => LPM_q_ivl_42645,
      b => LPM_q_ivl_42652,
      c => LPM_d0_ivl_42669,
      clk => clk,
      r => LPM_q_ivl_42659
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3291
  SboxInst_U129: not_masked
    port map (
      a => LPM_q_ivl_7105,
      b => LPM_d0_ivl_7107
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3349
  SboxInst_U13: not_masked
    port map (
      a => LPM_q_ivl_7627,
      b => LPM_d0_ivl_7629
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4885
  SboxInst_U130: and_HPC2
    port map (
      a => LPM_q_ivl_42617,
      b => LPM_q_ivl_42624,
      c => LPM_d0_ivl_42641,
      clk => clk,
      r => LPM_q_ivl_42631
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3290
  SboxInst_U131: not_masked
    port map (
      a => LPM_q_ivl_7096,
      b => LPM_d0_ivl_7098
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4884
  SboxInst_U132: and_HPC2
    port map (
      a => LPM_q_ivl_42589,
      b => LPM_q_ivl_42596,
      c => LPM_d0_ivl_42613,
      clk => clk,
      r => LPM_q_ivl_42603
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3289
  SboxInst_U133: not_masked
    port map (
      a => LPM_q_ivl_7087,
      b => LPM_d0_ivl_7089
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4883
  SboxInst_U134: and_HPC2
    port map (
      a => LPM_q_ivl_42561,
      b => LPM_q_ivl_42568,
      c => LPM_d0_ivl_42585,
      clk => clk,
      r => LPM_q_ivl_42575
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3288
  SboxInst_U135: not_masked
    port map (
      a => LPM_q_ivl_7078,
      b => LPM_d0_ivl_7080
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4882
  SboxInst_U136: and_HPC2
    port map (
      a => LPM_q_ivl_42533,
      b => LPM_q_ivl_42540,
      c => LPM_d0_ivl_42557,
      clk => clk,
      r => LPM_q_ivl_42547
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3287
  SboxInst_U137: not_masked
    port map (
      a => LPM_q_ivl_7069,
      b => LPM_d0_ivl_7071
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4881
  SboxInst_U138: and_HPC2
    port map (
      a => LPM_q_ivl_42505,
      b => LPM_q_ivl_42512,
      c => LPM_d0_ivl_42529,
      clk => clk,
      r => LPM_q_ivl_42519
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3286
  SboxInst_U139: not_masked
    port map (
      a => LPM_q_ivl_7060,
      b => LPM_d0_ivl_7062
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4943
  SboxInst_U14: and_HPC2
    port map (
      a => LPM_q_ivl_44279,
      b => LPM_q_ivl_44288,
      c => LPM_d0_ivl_44305,
      clk => clk,
      r => LPM_q_ivl_44295
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4880
  SboxInst_U140: and_HPC2
    port map (
      a => LPM_q_ivl_42477,
      b => LPM_q_ivl_42484,
      c => LPM_d0_ivl_42501,
      clk => clk,
      r => LPM_q_ivl_42491
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3285
  SboxInst_U141: not_masked
    port map (
      a => LPM_q_ivl_7051,
      b => LPM_d0_ivl_7053
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4879
  SboxInst_U142: and_HPC2
    port map (
      a => LPM_q_ivl_42449,
      b => LPM_q_ivl_42456,
      c => LPM_d0_ivl_42473,
      clk => clk,
      r => LPM_q_ivl_42463
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3284
  SboxInst_U143: not_masked
    port map (
      a => LPM_q_ivl_7042,
      b => LPM_d0_ivl_7044
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4878
  SboxInst_U144: and_HPC2
    port map (
      a => LPM_q_ivl_42421,
      b => LPM_q_ivl_42428,
      c => LPM_d0_ivl_42445,
      clk => clk,
      r => LPM_q_ivl_42435
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3283
  SboxInst_U145: not_masked
    port map (
      a => LPM_q_ivl_7033,
      b => LPM_d0_ivl_7035
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4877
  SboxInst_U146: and_HPC2
    port map (
      a => LPM_q_ivl_42393,
      b => LPM_q_ivl_42400,
      c => LPM_d0_ivl_42417,
      clk => clk,
      r => LPM_q_ivl_42407
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3282
  SboxInst_U147: not_masked
    port map (
      a => LPM_q_ivl_7024,
      b => LPM_d0_ivl_7026
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4876
  SboxInst_U148: and_HPC2
    port map (
      a => LPM_q_ivl_42365,
      b => LPM_q_ivl_42372,
      c => LPM_d0_ivl_42389,
      clk => clk,
      r => LPM_q_ivl_42379
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3281
  SboxInst_U149: not_masked
    port map (
      a => LPM_q_ivl_7015,
      b => LPM_d0_ivl_7017
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3348
  SboxInst_U15: not_masked
    port map (
      a => LPM_q_ivl_7618,
      b => LPM_d0_ivl_7620
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4875
  SboxInst_U150: and_HPC2
    port map (
      a => LPM_q_ivl_42337,
      b => LPM_q_ivl_42344,
      c => LPM_d0_ivl_42361,
      clk => clk,
      r => LPM_q_ivl_42351
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3280
  SboxInst_U151: not_masked
    port map (
      a => LPM_q_ivl_7006,
      b => LPM_d0_ivl_7008
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4874
  SboxInst_U152: and_HPC2
    port map (
      a => LPM_q_ivl_42309,
      b => LPM_q_ivl_42316,
      c => LPM_d0_ivl_42333,
      clk => clk,
      r => LPM_q_ivl_42323
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3279
  SboxInst_U153: not_masked
    port map (
      a => LPM_q_ivl_6997,
      b => LPM_d0_ivl_6999
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4873
  SboxInst_U154: and_HPC2
    port map (
      a => LPM_q_ivl_42281,
      b => LPM_q_ivl_42288,
      c => LPM_d0_ivl_42305,
      clk => clk,
      r => LPM_q_ivl_42295
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3278
  SboxInst_U155: not_masked
    port map (
      a => LPM_q_ivl_6988,
      b => LPM_d0_ivl_6990
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4872
  SboxInst_U156: and_HPC2
    port map (
      a => LPM_q_ivl_42253,
      b => LPM_q_ivl_42260,
      c => LPM_d0_ivl_42277,
      clk => clk,
      r => LPM_q_ivl_42267
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3277
  SboxInst_U157: not_masked
    port map (
      a => LPM_q_ivl_6979,
      b => LPM_d0_ivl_6981
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4871
  SboxInst_U158: and_HPC2
    port map (
      a => LPM_q_ivl_42223,
      b => LPM_q_ivl_42230,
      c => LPM_d0_ivl_42247,
      clk => clk,
      r => LPM_q_ivl_42237
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3276
  SboxInst_U159: not_masked
    port map (
      a => LPM_q_ivl_6970,
      b => LPM_d0_ivl_6972
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4942
  SboxInst_U16: and_HPC2
    port map (
      a => LPM_q_ivl_44249,
      b => LPM_q_ivl_44258,
      c => LPM_d0_ivl_44275,
      clk => clk,
      r => LPM_q_ivl_44265
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4870
  SboxInst_U160: and_HPC2
    port map (
      a => LPM_q_ivl_42195,
      b => LPM_q_ivl_42202,
      c => LPM_d0_ivl_42219,
      clk => clk,
      r => LPM_q_ivl_42209
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3275
  SboxInst_U161: not_masked
    port map (
      a => LPM_q_ivl_6961,
      b => LPM_d0_ivl_6963
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4869
  SboxInst_U162: and_HPC2
    port map (
      a => LPM_q_ivl_42165,
      b => LPM_q_ivl_42172,
      c => LPM_d0_ivl_42189,
      clk => clk,
      r => LPM_q_ivl_42179
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3274
  SboxInst_U163: not_masked
    port map (
      a => LPM_q_ivl_6952,
      b => LPM_d0_ivl_6954
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4868
  SboxInst_U164: and_HPC2
    port map (
      a => LPM_q_ivl_42137,
      b => LPM_q_ivl_42144,
      c => LPM_d0_ivl_42161,
      clk => clk,
      r => LPM_q_ivl_42151
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3273
  SboxInst_U165: not_masked
    port map (
      a => LPM_q_ivl_6943,
      b => LPM_d0_ivl_6945
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4867
  SboxInst_U166: and_HPC2
    port map (
      a => LPM_q_ivl_42109,
      b => LPM_q_ivl_42116,
      c => LPM_d0_ivl_42133,
      clk => clk,
      r => LPM_q_ivl_42123
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3272
  SboxInst_U167: not_masked
    port map (
      a => LPM_q_ivl_6934,
      b => LPM_d0_ivl_6936
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4866
  SboxInst_U168: and_HPC2
    port map (
      a => LPM_q_ivl_42081,
      b => LPM_q_ivl_42088,
      c => LPM_d0_ivl_42105,
      clk => clk,
      r => LPM_q_ivl_42095
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3271
  SboxInst_U169: not_masked
    port map (
      a => LPM_q_ivl_6925,
      b => LPM_d0_ivl_6927
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3347
  SboxInst_U17: not_masked
    port map (
      a => LPM_q_ivl_7609,
      b => LPM_d0_ivl_7611
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4865
  SboxInst_U170: and_HPC2
    port map (
      a => LPM_q_ivl_42053,
      b => LPM_q_ivl_42060,
      c => LPM_d0_ivl_42077,
      clk => clk,
      r => LPM_q_ivl_42067
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3270
  SboxInst_U171: not_masked
    port map (
      a => LPM_q_ivl_6916,
      b => LPM_d0_ivl_6918
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4864
  SboxInst_U172: and_HPC2
    port map (
      a => LPM_q_ivl_42025,
      b => LPM_q_ivl_42032,
      c => LPM_d0_ivl_42049,
      clk => clk,
      r => LPM_q_ivl_42039
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3269
  SboxInst_U173: not_masked
    port map (
      a => LPM_q_ivl_6907,
      b => LPM_d0_ivl_6909
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4863
  SboxInst_U174: and_HPC2
    port map (
      a => LPM_q_ivl_41997,
      b => LPM_q_ivl_42004,
      c => LPM_d0_ivl_42021,
      clk => clk,
      r => LPM_q_ivl_42011
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3268
  SboxInst_U175: not_masked
    port map (
      a => LPM_q_ivl_6898,
      b => LPM_d0_ivl_6900
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4862
  SboxInst_U176: and_HPC2
    port map (
      a => LPM_q_ivl_41969,
      b => LPM_q_ivl_41976,
      c => LPM_d0_ivl_41993,
      clk => clk,
      r => LPM_q_ivl_41983
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3267
  SboxInst_U177: not_masked
    port map (
      a => LPM_q_ivl_6889,
      b => LPM_d0_ivl_6891
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4861
  SboxInst_U178: and_HPC2
    port map (
      a => LPM_q_ivl_41941,
      b => LPM_q_ivl_41948,
      c => LPM_d0_ivl_41965,
      clk => clk,
      r => LPM_q_ivl_41955
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3266
  SboxInst_U179: not_masked
    port map (
      a => LPM_q_ivl_6880,
      b => LPM_d0_ivl_6882
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4941
  SboxInst_U18: and_HPC2
    port map (
      a => LPM_q_ivl_44219,
      b => LPM_q_ivl_44228,
      c => LPM_d0_ivl_44245,
      clk => clk,
      r => LPM_q_ivl_44235
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4860
  SboxInst_U180: and_HPC2
    port map (
      a => LPM_q_ivl_41913,
      b => LPM_q_ivl_41920,
      c => LPM_d0_ivl_41937,
      clk => clk,
      r => LPM_q_ivl_41927
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3265
  SboxInst_U181: not_masked
    port map (
      a => LPM_q_ivl_6871,
      b => LPM_d0_ivl_6873
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4859
  SboxInst_U182: and_HPC2
    port map (
      a => LPM_q_ivl_41883,
      b => LPM_q_ivl_41892,
      c => LPM_d0_ivl_41909,
      clk => clk,
      r => LPM_q_ivl_41899
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3264
  SboxInst_U183: not_masked
    port map (
      a => LPM_q_ivl_6862,
      b => LPM_d0_ivl_6864
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4858
  SboxInst_U184: and_HPC2
    port map (
      a => LPM_q_ivl_41853,
      b => LPM_q_ivl_41862,
      c => LPM_d0_ivl_41879,
      clk => clk,
      r => LPM_q_ivl_41869
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3263
  SboxInst_U185: not_masked
    port map (
      a => LPM_q_ivl_6853,
      b => LPM_d0_ivl_6855
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4857
  SboxInst_U186: and_HPC2
    port map (
      a => LPM_q_ivl_41823,
      b => LPM_q_ivl_41832,
      c => LPM_d0_ivl_41849,
      clk => clk,
      r => LPM_q_ivl_41839
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3262
  SboxInst_U187: not_masked
    port map (
      a => LPM_q_ivl_6844,
      b => LPM_d0_ivl_6846
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4856
  SboxInst_U188: and_HPC2
    port map (
      a => LPM_q_ivl_41793,
      b => LPM_q_ivl_41802,
      c => LPM_d0_ivl_41819,
      clk => clk,
      r => LPM_q_ivl_41809
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3261
  SboxInst_U189: not_masked
    port map (
      a => LPM_q_ivl_6835,
      b => LPM_d0_ivl_6837
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3346
  SboxInst_U19: not_masked
    port map (
      a => LPM_q_ivl_7600,
      b => LPM_d0_ivl_7602
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4855
  SboxInst_U190: and_HPC2
    port map (
      a => LPM_q_ivl_41763,
      b => LPM_q_ivl_41772,
      c => LPM_d0_ivl_41789,
      clk => clk,
      r => LPM_q_ivl_41779
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3260
  SboxInst_U191: not_masked
    port map (
      a => LPM_q_ivl_6826,
      b => LPM_d0_ivl_6828
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4854
  SboxInst_U192: and_HPC2
    port map (
      a => LPM_q_ivl_41733,
      b => LPM_q_ivl_41742,
      c => LPM_d0_ivl_41759,
      clk => clk,
      r => LPM_q_ivl_41749
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3259
  SboxInst_U193: not_masked
    port map (
      a => LPM_q_ivl_6817,
      b => LPM_d0_ivl_6819
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4853
  SboxInst_U194: and_HPC2
    port map (
      a => LPM_q_ivl_41703,
      b => LPM_q_ivl_41712,
      c => LPM_d0_ivl_41729,
      clk => clk,
      r => LPM_q_ivl_41719
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3258
  SboxInst_U195: not_masked
    port map (
      a => LPM_q_ivl_6808,
      b => LPM_d0_ivl_6810
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4852
  SboxInst_U196: and_HPC2
    port map (
      a => LPM_q_ivl_41673,
      b => LPM_q_ivl_41682,
      c => LPM_d0_ivl_41699,
      clk => clk,
      r => LPM_q_ivl_41689
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3257
  SboxInst_U197: not_masked
    port map (
      a => LPM_q_ivl_6799,
      b => LPM_d0_ivl_6801
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4851
  SboxInst_U198: and_HPC2
    port map (
      a => LPM_q_ivl_41643,
      b => LPM_q_ivl_41652,
      c => LPM_d0_ivl_41669,
      clk => clk,
      r => LPM_q_ivl_41659
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3256
  SboxInst_U199: not_masked
    port map (
      a => LPM_q_ivl_6790,
      b => LPM_d0_ivl_6792
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4949
  SboxInst_U2: and_HPC2
    port map (
      a => LPM_q_ivl_44459,
      b => LPM_q_ivl_44468,
      c => LPM_d0_ivl_44485,
      clk => clk,
      r => LPM_q_ivl_44475
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4940
  SboxInst_U20: and_HPC2
    port map (
      a => LPM_q_ivl_44189,
      b => LPM_q_ivl_44198,
      c => LPM_d0_ivl_44215,
      clk => clk,
      r => LPM_q_ivl_44205
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4850
  SboxInst_U200: and_HPC2
    port map (
      a => LPM_q_ivl_41613,
      b => LPM_q_ivl_41622,
      c => LPM_d0_ivl_41639,
      clk => clk,
      r => LPM_q_ivl_41629
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3255
  SboxInst_U201: not_masked
    port map (
      a => LPM_q_ivl_6781,
      b => LPM_d0_ivl_6783
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4849
  SboxInst_U202: and_HPC2
    port map (
      a => LPM_q_ivl_41583,
      b => LPM_q_ivl_41592,
      c => LPM_d0_ivl_41609,
      clk => clk,
      r => LPM_q_ivl_41599
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3254
  SboxInst_U203: not_masked
    port map (
      a => LPM_q_ivl_6772,
      b => LPM_d0_ivl_6774
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4848
  SboxInst_U204: and_HPC2
    port map (
      a => LPM_q_ivl_41553,
      b => LPM_q_ivl_41562,
      c => LPM_d0_ivl_41579,
      clk => clk,
      r => LPM_q_ivl_41569
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3253
  SboxInst_U205: not_masked
    port map (
      a => LPM_q_ivl_6763,
      b => LPM_d0_ivl_6765
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4847
  SboxInst_U206: and_HPC2
    port map (
      a => LPM_q_ivl_41523,
      b => LPM_q_ivl_41532,
      c => LPM_d0_ivl_41549,
      clk => clk,
      r => LPM_q_ivl_41539
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3252
  SboxInst_U207: not_masked
    port map (
      a => LPM_q_ivl_6754,
      b => LPM_d0_ivl_6756
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4846
  SboxInst_U208: and_HPC2
    port map (
      a => LPM_q_ivl_41493,
      b => LPM_q_ivl_41502,
      c => LPM_d0_ivl_41519,
      clk => clk,
      r => LPM_q_ivl_41509
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3251
  SboxInst_U209: not_masked
    port map (
      a => LPM_q_ivl_6745,
      b => LPM_d0_ivl_6747
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3345
  SboxInst_U21: not_masked
    port map (
      a => LPM_q_ivl_7591,
      b => LPM_d0_ivl_7593
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4845
  SboxInst_U210: and_HPC2
    port map (
      a => LPM_q_ivl_41463,
      b => LPM_q_ivl_41472,
      c => LPM_d0_ivl_41489,
      clk => clk,
      r => LPM_q_ivl_41479
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3250
  SboxInst_U211: not_masked
    port map (
      a => LPM_q_ivl_6736,
      b => LPM_d0_ivl_6738
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4844
  SboxInst_U212: and_HPC2
    port map (
      a => LPM_q_ivl_41433,
      b => LPM_q_ivl_41442,
      c => LPM_d0_ivl_41459,
      clk => clk,
      r => LPM_q_ivl_41449
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3249
  SboxInst_U213: not_masked
    port map (
      a => LPM_q_ivl_6727,
      b => LPM_d0_ivl_6729
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4843
  SboxInst_U214: and_HPC2
    port map (
      a => LPM_q_ivl_41403,
      b => LPM_q_ivl_41412,
      c => LPM_d0_ivl_41429,
      clk => clk,
      r => LPM_q_ivl_41419
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3248
  SboxInst_U215: not_masked
    port map (
      a => LPM_q_ivl_6718,
      b => LPM_d0_ivl_6720
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4842
  SboxInst_U216: and_HPC2
    port map (
      a => LPM_q_ivl_41373,
      b => LPM_q_ivl_41382,
      c => LPM_d0_ivl_41399,
      clk => clk,
      r => LPM_q_ivl_41389
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3247
  SboxInst_U217: not_masked
    port map (
      a => LPM_q_ivl_6709,
      b => LPM_d0_ivl_6711
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4841
  SboxInst_U218: and_HPC2
    port map (
      a => LPM_q_ivl_41343,
      b => LPM_q_ivl_41352,
      c => LPM_d0_ivl_41369,
      clk => clk,
      r => LPM_q_ivl_41359
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3246
  SboxInst_U219: not_masked
    port map (
      a => LPM_q_ivl_6700,
      b => LPM_d0_ivl_6702
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4939
  SboxInst_U22: and_HPC2
    port map (
      a => LPM_q_ivl_44159,
      b => LPM_q_ivl_44168,
      c => LPM_d0_ivl_44185,
      clk => clk,
      r => LPM_q_ivl_44175
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4840
  SboxInst_U220: and_HPC2
    port map (
      a => LPM_q_ivl_41313,
      b => LPM_q_ivl_41322,
      c => LPM_d0_ivl_41339,
      clk => clk,
      r => LPM_q_ivl_41329
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3245
  SboxInst_U221: not_masked
    port map (
      a => LPM_q_ivl_6691,
      b => LPM_d0_ivl_6693
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4839
  SboxInst_U222: and_HPC2
    port map (
      a => LPM_q_ivl_41283,
      b => LPM_q_ivl_41292,
      c => LPM_d0_ivl_41309,
      clk => clk,
      r => LPM_q_ivl_41299
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3244
  SboxInst_U223: not_masked
    port map (
      a => LPM_q_ivl_6682,
      b => LPM_d0_ivl_6684
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4838
  SboxInst_U224: and_HPC2
    port map (
      a => LPM_q_ivl_41253,
      b => LPM_q_ivl_41262,
      c => LPM_d0_ivl_41279,
      clk => clk,
      r => LPM_q_ivl_41269
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3243
  SboxInst_U225: not_masked
    port map (
      a => LPM_q_ivl_6673,
      b => LPM_d0_ivl_6675
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4837
  SboxInst_U226: and_HPC2
    port map (
      a => LPM_q_ivl_41223,
      b => LPM_q_ivl_41232,
      c => LPM_d0_ivl_41249,
      clk => clk,
      r => LPM_q_ivl_41239
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3242
  SboxInst_U227: not_masked
    port map (
      a => LPM_q_ivl_6664,
      b => LPM_d0_ivl_6666
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4836
  SboxInst_U228: and_HPC2
    port map (
      a => LPM_q_ivl_41193,
      b => LPM_q_ivl_41202,
      c => LPM_d0_ivl_41219,
      clk => clk,
      r => LPM_q_ivl_41209
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3241
  SboxInst_U229: not_masked
    port map (
      a => LPM_q_ivl_6655,
      b => LPM_d0_ivl_6657
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3344
  SboxInst_U23: not_masked
    port map (
      a => LPM_q_ivl_7582,
      b => LPM_d0_ivl_7584
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4835
  SboxInst_U230: and_HPC2
    port map (
      a => LPM_q_ivl_41163,
      b => LPM_q_ivl_41172,
      c => LPM_d0_ivl_41189,
      clk => clk,
      r => LPM_q_ivl_41179
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3240
  SboxInst_U231: not_masked
    port map (
      a => LPM_q_ivl_6646,
      b => LPM_d0_ivl_6648
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4834
  SboxInst_U232: and_HPC2
    port map (
      a => LPM_q_ivl_41133,
      b => LPM_q_ivl_41142,
      c => LPM_d0_ivl_41159,
      clk => clk,
      r => LPM_q_ivl_41149
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3239
  SboxInst_U233: not_masked
    port map (
      a => LPM_q_ivl_6637,
      b => LPM_d0_ivl_6639
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4833
  SboxInst_U234: and_HPC2
    port map (
      a => LPM_q_ivl_41103,
      b => LPM_q_ivl_41112,
      c => LPM_d0_ivl_41129,
      clk => clk,
      r => LPM_q_ivl_41119
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3238
  SboxInst_U235: not_masked
    port map (
      a => LPM_q_ivl_6628,
      b => LPM_d0_ivl_6630
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4832
  SboxInst_U236: and_HPC2
    port map (
      a => LPM_q_ivl_41073,
      b => LPM_q_ivl_41082,
      c => LPM_d0_ivl_41099,
      clk => clk,
      r => LPM_q_ivl_41089
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3237
  SboxInst_U237: not_masked
    port map (
      a => LPM_q_ivl_6619,
      b => LPM_d0_ivl_6621
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4831
  SboxInst_U238: and_HPC2
    port map (
      a => LPM_q_ivl_41043,
      b => LPM_q_ivl_41052,
      c => LPM_d0_ivl_41069,
      clk => clk,
      r => LPM_q_ivl_41059
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3236
  SboxInst_U239: not_masked
    port map (
      a => LPM_q_ivl_6610,
      b => LPM_d0_ivl_6612
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4938
  SboxInst_U24: and_HPC2
    port map (
      a => LPM_q_ivl_44129,
      b => LPM_q_ivl_44138,
      c => LPM_d0_ivl_44155,
      clk => clk,
      r => LPM_q_ivl_44145
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4830
  SboxInst_U240: and_HPC2
    port map (
      a => LPM_q_ivl_41013,
      b => LPM_q_ivl_41022,
      c => LPM_d0_ivl_41039,
      clk => clk,
      r => LPM_q_ivl_41029
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3235
  SboxInst_U241: not_masked
    port map (
      a => LPM_q_ivl_6601,
      b => LPM_d0_ivl_6603
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4829
  SboxInst_U242: and_HPC2
    port map (
      a => LPM_q_ivl_40983,
      b => LPM_q_ivl_40992,
      c => LPM_d0_ivl_41009,
      clk => clk,
      r => LPM_q_ivl_40999
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3234
  SboxInst_U243: not_masked
    port map (
      a => LPM_q_ivl_6592,
      b => LPM_d0_ivl_6594
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4828
  SboxInst_U244: and_HPC2
    port map (
      a => LPM_q_ivl_40953,
      b => LPM_q_ivl_40962,
      c => LPM_d0_ivl_40979,
      clk => clk,
      r => LPM_q_ivl_40969
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3233
  SboxInst_U245: not_masked
    port map (
      a => LPM_q_ivl_6583,
      b => LPM_d0_ivl_6585
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4827
  SboxInst_U246: and_HPC2
    port map (
      a => LPM_q_ivl_40923,
      b => LPM_q_ivl_40932,
      c => LPM_d0_ivl_40949,
      clk => clk,
      r => LPM_q_ivl_40939
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3232
  SboxInst_U247: not_masked
    port map (
      a => LPM_q_ivl_6574,
      b => LPM_d0_ivl_6576
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4826
  SboxInst_U248: and_HPC2
    port map (
      a => LPM_q_ivl_40893,
      b => LPM_q_ivl_40902,
      c => LPM_d0_ivl_40919,
      clk => clk,
      r => LPM_q_ivl_40909
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3231
  SboxInst_U249: not_masked
    port map (
      a => LPM_q_ivl_6565,
      b => LPM_d0_ivl_6567
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3343
  SboxInst_U25: not_masked
    port map (
      a => LPM_q_ivl_7573,
      b => LPM_d0_ivl_7575
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4825
  SboxInst_U250: and_HPC2
    port map (
      a => LPM_q_ivl_40863,
      b => LPM_q_ivl_40872,
      c => LPM_d0_ivl_40889,
      clk => clk,
      r => LPM_q_ivl_40879
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3230
  SboxInst_U251: not_masked
    port map (
      a => LPM_q_ivl_6556,
      b => LPM_d0_ivl_6558
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4824
  SboxInst_U252: and_HPC2
    port map (
      a => LPM_q_ivl_40833,
      b => LPM_q_ivl_40842,
      c => LPM_d0_ivl_40859,
      clk => clk,
      r => LPM_q_ivl_40849
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3229
  SboxInst_U253: not_masked
    port map (
      a => LPM_q_ivl_6547,
      b => LPM_d0_ivl_6549
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4823
  SboxInst_U254: and_HPC2
    port map (
      a => LPM_q_ivl_40803,
      b => LPM_q_ivl_40812,
      c => LPM_d0_ivl_40829,
      clk => clk,
      r => LPM_q_ivl_40819
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3228
  SboxInst_U255: not_masked
    port map (
      a => LPM_q_ivl_6538,
      b => LPM_d0_ivl_6540
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4822
  SboxInst_U256: and_HPC2
    port map (
      a => LPM_q_ivl_40773,
      b => LPM_q_ivl_40782,
      c => LPM_d0_ivl_40799,
      clk => clk,
      r => LPM_q_ivl_40789
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4821
  SboxInst_U257: nor_HPC2
    port map (
      a => LPM_q_ivl_40745,
      b => LPM_q_ivl_40752,
      c => LPM_d0_ivl_40769,
      clk => clk,
      r => LPM_q_ivl_40759
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4820
  SboxInst_U258: nor_HPC2
    port map (
      a => LPM_q_ivl_40715,
      b => LPM_q_ivl_40722,
      c => LPM_d0_ivl_40739,
      clk => clk,
      r => LPM_q_ivl_40729
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4819
  SboxInst_U259: nor_HPC2
    port map (
      a => LPM_q_ivl_40685,
      b => LPM_q_ivl_40692,
      c => LPM_d0_ivl_40709,
      clk => clk,
      r => LPM_q_ivl_40699
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4937
  SboxInst_U26: and_HPC2
    port map (
      a => LPM_q_ivl_44099,
      b => LPM_q_ivl_44108,
      c => LPM_d0_ivl_44125,
      clk => clk,
      r => LPM_q_ivl_44115
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4818
  SboxInst_U260: nor_HPC2
    port map (
      a => LPM_q_ivl_40655,
      b => LPM_q_ivl_40662,
      c => LPM_d0_ivl_40679,
      clk => clk,
      r => LPM_q_ivl_40669
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4817
  SboxInst_U261: nor_HPC2
    port map (
      a => LPM_q_ivl_40625,
      b => LPM_q_ivl_40632,
      c => LPM_d0_ivl_40649,
      clk => clk,
      r => LPM_q_ivl_40639
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4816
  SboxInst_U262: nor_HPC2
    port map (
      a => LPM_q_ivl_40595,
      b => LPM_q_ivl_40602,
      c => LPM_d0_ivl_40619,
      clk => clk,
      r => LPM_q_ivl_40609
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4815
  SboxInst_U263: nor_HPC2
    port map (
      a => LPM_q_ivl_40565,
      b => LPM_q_ivl_40572,
      c => LPM_d0_ivl_40589,
      clk => clk,
      r => LPM_q_ivl_40579
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4814
  SboxInst_U264: nor_HPC2
    port map (
      a => LPM_q_ivl_40535,
      b => LPM_q_ivl_40542,
      c => LPM_d0_ivl_40559,
      clk => clk,
      r => LPM_q_ivl_40549
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4813
  SboxInst_U265: nor_HPC2
    port map (
      a => LPM_q_ivl_40505,
      b => LPM_q_ivl_40512,
      c => LPM_d0_ivl_40529,
      clk => clk,
      r => LPM_q_ivl_40519
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4812
  SboxInst_U266: nor_HPC2
    port map (
      a => LPM_q_ivl_40475,
      b => LPM_q_ivl_40482,
      c => LPM_d0_ivl_40499,
      clk => clk,
      r => LPM_q_ivl_40489
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4811
  SboxInst_U267: nor_HPC2
    port map (
      a => LPM_q_ivl_40445,
      b => LPM_q_ivl_40452,
      c => LPM_d0_ivl_40469,
      clk => clk,
      r => LPM_q_ivl_40459
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4810
  SboxInst_U268: nor_HPC2
    port map (
      a => LPM_q_ivl_40415,
      b => LPM_q_ivl_40422,
      c => LPM_d0_ivl_40439,
      clk => clk,
      r => LPM_q_ivl_40429
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4809
  SboxInst_U269: nor_HPC2
    port map (
      a => LPM_q_ivl_40385,
      b => LPM_q_ivl_40392,
      c => LPM_d0_ivl_40409,
      clk => clk,
      r => LPM_q_ivl_40399
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3342
  SboxInst_U27: not_masked
    port map (
      a => LPM_q_ivl_7564,
      b => LPM_d0_ivl_7566
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4808
  SboxInst_U270: nor_HPC2
    port map (
      a => LPM_q_ivl_40355,
      b => LPM_q_ivl_40362,
      c => LPM_d0_ivl_40379,
      clk => clk,
      r => LPM_q_ivl_40369
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4807
  SboxInst_U271: nor_HPC2
    port map (
      a => LPM_q_ivl_40325,
      b => LPM_q_ivl_40332,
      c => LPM_d0_ivl_40349,
      clk => clk,
      r => LPM_q_ivl_40339
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4806
  SboxInst_U272: nor_HPC2
    port map (
      a => LPM_q_ivl_40295,
      b => LPM_q_ivl_40302,
      c => LPM_d0_ivl_40319,
      clk => clk,
      r => LPM_q_ivl_40309
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4805
  SboxInst_U273: nor_HPC2
    port map (
      a => LPM_q_ivl_40265,
      b => LPM_q_ivl_40272,
      c => LPM_d0_ivl_40289,
      clk => clk,
      r => LPM_q_ivl_40279
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4804
  SboxInst_U274: nor_HPC2
    port map (
      a => LPM_q_ivl_40235,
      b => LPM_q_ivl_40242,
      c => LPM_d0_ivl_40259,
      clk => clk,
      r => LPM_q_ivl_40249
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4803
  SboxInst_U275: nor_HPC2
    port map (
      a => LPM_q_ivl_40205,
      b => LPM_q_ivl_40212,
      c => LPM_d0_ivl_40229,
      clk => clk,
      r => LPM_q_ivl_40219
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4802
  SboxInst_U276: nor_HPC2
    port map (
      a => LPM_q_ivl_40175,
      b => LPM_q_ivl_40182,
      c => LPM_d0_ivl_40199,
      clk => clk,
      r => LPM_q_ivl_40189
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4801
  SboxInst_U277: nor_HPC2
    port map (
      a => LPM_q_ivl_40145,
      b => LPM_q_ivl_40152,
      c => LPM_d0_ivl_40169,
      clk => clk,
      r => LPM_q_ivl_40159
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4800
  SboxInst_U278: nor_HPC2
    port map (
      a => LPM_q_ivl_40115,
      b => LPM_q_ivl_40122,
      c => LPM_d0_ivl_40139,
      clk => clk,
      r => LPM_q_ivl_40129
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4799
  SboxInst_U279: nor_HPC2
    port map (
      a => LPM_q_ivl_40085,
      b => LPM_q_ivl_40092,
      c => LPM_d0_ivl_40109,
      clk => clk,
      r => LPM_q_ivl_40099
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4936
  SboxInst_U28: and_HPC2
    port map (
      a => LPM_q_ivl_44069,
      b => LPM_q_ivl_44078,
      c => LPM_d0_ivl_44095,
      clk => clk,
      r => LPM_q_ivl_44085
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4798
  SboxInst_U280: nor_HPC2
    port map (
      a => LPM_q_ivl_40055,
      b => LPM_q_ivl_40062,
      c => LPM_d0_ivl_40079,
      clk => clk,
      r => LPM_q_ivl_40069
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4797
  SboxInst_U281: nor_HPC2
    port map (
      a => LPM_q_ivl_40025,
      b => LPM_q_ivl_40032,
      c => LPM_d0_ivl_40049,
      clk => clk,
      r => LPM_q_ivl_40039
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4796
  SboxInst_U282: nor_HPC2
    port map (
      a => LPM_q_ivl_39995,
      b => LPM_q_ivl_40002,
      c => LPM_d0_ivl_40019,
      clk => clk,
      r => LPM_q_ivl_40009
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4795
  SboxInst_U283: nor_HPC2
    port map (
      a => LPM_q_ivl_39965,
      b => LPM_q_ivl_39972,
      c => LPM_d0_ivl_39989,
      clk => clk,
      r => LPM_q_ivl_39979
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4794
  SboxInst_U284: nor_HPC2
    port map (
      a => LPM_q_ivl_39935,
      b => LPM_q_ivl_39942,
      c => LPM_d0_ivl_39959,
      clk => clk,
      r => LPM_q_ivl_39949
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4793
  SboxInst_U285: nor_HPC2
    port map (
      a => LPM_q_ivl_39905,
      b => LPM_q_ivl_39912,
      c => LPM_d0_ivl_39929,
      clk => clk,
      r => LPM_q_ivl_39919
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4792
  SboxInst_U286: nor_HPC2
    port map (
      a => LPM_q_ivl_39875,
      b => LPM_q_ivl_39882,
      c => LPM_d0_ivl_39899,
      clk => clk,
      r => LPM_q_ivl_39889
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4791
  SboxInst_U287: nor_HPC2
    port map (
      a => LPM_q_ivl_39845,
      b => LPM_q_ivl_39852,
      c => LPM_d0_ivl_39869,
      clk => clk,
      r => LPM_q_ivl_39859
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4790
  SboxInst_U288: nor_HPC2
    port map (
      a => LPM_q_ivl_39815,
      b => LPM_q_ivl_39822,
      c => LPM_d0_ivl_39839,
      clk => clk,
      r => LPM_q_ivl_39829
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4789
  SboxInst_U289: nor_HPC2
    port map (
      a => LPM_q_ivl_39785,
      b => LPM_q_ivl_39792,
      c => LPM_d0_ivl_39809,
      clk => clk,
      r => LPM_q_ivl_39799
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3341
  SboxInst_U29: not_masked
    port map (
      a => LPM_q_ivl_7555,
      b => LPM_d0_ivl_7557
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4788
  SboxInst_U290: nor_HPC2
    port map (
      a => LPM_q_ivl_39755,
      b => LPM_q_ivl_39762,
      c => LPM_d0_ivl_39779,
      clk => clk,
      r => LPM_q_ivl_39769
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4787
  SboxInst_U291: nor_HPC2
    port map (
      a => LPM_q_ivl_39725,
      b => LPM_q_ivl_39732,
      c => LPM_d0_ivl_39749,
      clk => clk,
      r => LPM_q_ivl_39739
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4786
  SboxInst_U292: nor_HPC2
    port map (
      a => LPM_q_ivl_39695,
      b => LPM_q_ivl_39702,
      c => LPM_d0_ivl_39719,
      clk => clk,
      r => LPM_q_ivl_39709
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4785
  SboxInst_U293: nor_HPC2
    port map (
      a => LPM_q_ivl_39665,
      b => LPM_q_ivl_39672,
      c => LPM_d0_ivl_39689,
      clk => clk,
      r => LPM_q_ivl_39679
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4784
  SboxInst_U294: nor_HPC2
    port map (
      a => LPM_q_ivl_39635,
      b => LPM_q_ivl_39642,
      c => LPM_d0_ivl_39659,
      clk => clk,
      r => LPM_q_ivl_39649
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4783
  SboxInst_U295: nor_HPC2
    port map (
      a => LPM_q_ivl_39605,
      b => LPM_q_ivl_39612,
      c => LPM_d0_ivl_39629,
      clk => clk,
      r => LPM_q_ivl_39619
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4782
  SboxInst_U296: nor_HPC2
    port map (
      a => LPM_q_ivl_39575,
      b => LPM_q_ivl_39582,
      c => LPM_d0_ivl_39599,
      clk => clk,
      r => LPM_q_ivl_39589
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4781
  SboxInst_U297: nor_HPC2
    port map (
      a => LPM_q_ivl_39545,
      b => LPM_q_ivl_39552,
      c => LPM_d0_ivl_39569,
      clk => clk,
      r => LPM_q_ivl_39559
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4780
  SboxInst_U298: nor_HPC2
    port map (
      a => LPM_q_ivl_39515,
      b => LPM_q_ivl_39522,
      c => LPM_d0_ivl_39539,
      clk => clk,
      r => LPM_q_ivl_39529
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4779
  SboxInst_U299: nor_HPC2
    port map (
      a => LPM_q_ivl_39485,
      b => LPM_q_ivl_39492,
      c => LPM_d0_ivl_39509,
      clk => clk,
      r => LPM_q_ivl_39499
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3354
  SboxInst_U3: not_masked
    port map (
      a => LPM_q_ivl_7672,
      b => LPM_d0_ivl_7674
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4935
  SboxInst_U30: and_HPC2
    port map (
      a => LPM_q_ivl_44039,
      b => LPM_q_ivl_44048,
      c => LPM_d0_ivl_44065,
      clk => clk,
      r => LPM_q_ivl_44055
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4778
  SboxInst_U300: nor_HPC2
    port map (
      a => LPM_q_ivl_39455,
      b => LPM_q_ivl_39462,
      c => LPM_d0_ivl_39479,
      clk => clk,
      r => LPM_q_ivl_39469
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4777
  SboxInst_U301: nor_HPC2
    port map (
      a => LPM_q_ivl_39425,
      b => LPM_q_ivl_39432,
      c => LPM_d0_ivl_39449,
      clk => clk,
      r => LPM_q_ivl_39439
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4776
  SboxInst_U302: nor_HPC2
    port map (
      a => LPM_q_ivl_39395,
      b => LPM_q_ivl_39402,
      c => LPM_d0_ivl_39419,
      clk => clk,
      r => LPM_q_ivl_39409
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4775
  SboxInst_U303: nor_HPC2
    port map (
      a => LPM_q_ivl_39365,
      b => LPM_q_ivl_39372,
      c => LPM_d0_ivl_39389,
      clk => clk,
      r => LPM_q_ivl_39379
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4774
  SboxInst_U304: nor_HPC2
    port map (
      a => LPM_q_ivl_39335,
      b => LPM_q_ivl_39342,
      c => LPM_d0_ivl_39359,
      clk => clk,
      r => LPM_q_ivl_39349
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4773
  SboxInst_U305: nor_HPC2
    port map (
      a => LPM_q_ivl_39305,
      b => LPM_q_ivl_39312,
      c => LPM_d0_ivl_39329,
      clk => clk,
      r => LPM_q_ivl_39319
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4772
  SboxInst_U306: nor_HPC2
    port map (
      a => LPM_q_ivl_39275,
      b => LPM_q_ivl_39282,
      c => LPM_d0_ivl_39299,
      clk => clk,
      r => LPM_q_ivl_39289
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4771
  SboxInst_U307: nor_HPC2
    port map (
      a => LPM_q_ivl_39245,
      b => LPM_q_ivl_39252,
      c => LPM_d0_ivl_39269,
      clk => clk,
      r => LPM_q_ivl_39259
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4770
  SboxInst_U308: nor_HPC2
    port map (
      a => LPM_q_ivl_39215,
      b => LPM_q_ivl_39222,
      c => LPM_d0_ivl_39239,
      clk => clk,
      r => LPM_q_ivl_39229
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4769
  SboxInst_U309: nor_HPC2
    port map (
      a => LPM_q_ivl_39185,
      b => LPM_q_ivl_39192,
      c => LPM_d0_ivl_39209,
      clk => clk,
      r => LPM_q_ivl_39199
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3340
  SboxInst_U31: not_masked
    port map (
      a => LPM_q_ivl_7546,
      b => LPM_d0_ivl_7548
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4768
  SboxInst_U310: nor_HPC2
    port map (
      a => LPM_q_ivl_39155,
      b => LPM_q_ivl_39162,
      c => LPM_d0_ivl_39179,
      clk => clk,
      r => LPM_q_ivl_39169
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4767
  SboxInst_U311: nor_HPC2
    port map (
      a => LPM_q_ivl_39125,
      b => LPM_q_ivl_39132,
      c => LPM_d0_ivl_39149,
      clk => clk,
      r => LPM_q_ivl_39139
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4766
  SboxInst_U312: nor_HPC2
    port map (
      a => LPM_q_ivl_39095,
      b => LPM_q_ivl_39102,
      c => LPM_d0_ivl_39119,
      clk => clk,
      r => LPM_q_ivl_39109
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4765
  SboxInst_U313: nor_HPC2
    port map (
      a => LPM_q_ivl_39065,
      b => LPM_q_ivl_39072,
      c => LPM_d0_ivl_39089,
      clk => clk,
      r => LPM_q_ivl_39079
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4764
  SboxInst_U314: nor_HPC2
    port map (
      a => LPM_q_ivl_39035,
      b => LPM_q_ivl_39042,
      c => LPM_d0_ivl_39059,
      clk => clk,
      r => LPM_q_ivl_39049
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4763
  SboxInst_U315: nor_HPC2
    port map (
      a => LPM_q_ivl_39005,
      b => LPM_q_ivl_39012,
      c => LPM_d0_ivl_39029,
      clk => clk,
      r => LPM_q_ivl_39019
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4762
  SboxInst_U316: nor_HPC2
    port map (
      a => LPM_q_ivl_38975,
      b => LPM_q_ivl_38982,
      c => LPM_d0_ivl_38999,
      clk => clk,
      r => LPM_q_ivl_38989
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4761
  SboxInst_U317: nor_HPC2
    port map (
      a => LPM_q_ivl_38945,
      b => LPM_q_ivl_38952,
      c => LPM_d0_ivl_38969,
      clk => clk,
      r => LPM_q_ivl_38959
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4760
  SboxInst_U318: nor_HPC2
    port map (
      a => LPM_q_ivl_38915,
      b => LPM_q_ivl_38922,
      c => LPM_d0_ivl_38939,
      clk => clk,
      r => LPM_q_ivl_38929
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4759
  SboxInst_U319: nor_HPC2
    port map (
      a => LPM_q_ivl_38885,
      b => LPM_q_ivl_38892,
      c => LPM_d0_ivl_38909,
      clk => clk,
      r => LPM_q_ivl_38899
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4934
  SboxInst_U32: and_HPC2
    port map (
      a => LPM_q_ivl_44009,
      b => LPM_q_ivl_44018,
      c => LPM_d0_ivl_44035,
      clk => clk,
      r => LPM_q_ivl_44025
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4758
  SboxInst_U320: nor_HPC2
    port map (
      a => LPM_q_ivl_38855,
      b => LPM_q_ivl_38862,
      c => LPM_d0_ivl_38879,
      clk => clk,
      r => LPM_q_ivl_38869
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3227
  SboxInst_U321: not_masked
    port map (
      a => LPM_q_ivl_6529,
      b => LPM_d0_ivl_6531
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4757
  SboxInst_U322: nor_HPC2
    port map (
      a => LPM_q_ivl_38825,
      b => LPM_q_ivl_38832,
      c => LPM_d0_ivl_38849,
      clk => clk,
      r => LPM_q_ivl_38839
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3226
  SboxInst_U323: not_masked
    port map (
      a => LPM_q_ivl_6522,
      b => LPM_d0_ivl_6524
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4756
  SboxInst_U324: nor_HPC2
    port map (
      a => LPM_q_ivl_38795,
      b => LPM_q_ivl_38802,
      c => LPM_d0_ivl_38819,
      clk => clk,
      r => LPM_q_ivl_38809
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3225
  SboxInst_U325: not_masked
    port map (
      a => LPM_q_ivl_6515,
      b => LPM_d0_ivl_6517
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4755
  SboxInst_U326: nor_HPC2
    port map (
      a => LPM_q_ivl_38765,
      b => LPM_q_ivl_38772,
      c => LPM_d0_ivl_38789,
      clk => clk,
      r => LPM_q_ivl_38779
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3224
  SboxInst_U327: not_masked
    port map (
      a => LPM_q_ivl_6508,
      b => LPM_d0_ivl_6510
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4754
  SboxInst_U328: nor_HPC2
    port map (
      a => LPM_q_ivl_38735,
      b => LPM_q_ivl_38742,
      c => LPM_d0_ivl_38759,
      clk => clk,
      r => LPM_q_ivl_38749
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3223
  SboxInst_U329: not_masked
    port map (
      a => LPM_q_ivl_6501,
      b => LPM_d0_ivl_6503
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3339
  SboxInst_U33: not_masked
    port map (
      a => LPM_q_ivl_7537,
      b => LPM_d0_ivl_7539
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4753
  SboxInst_U330: nor_HPC2
    port map (
      a => LPM_q_ivl_38705,
      b => LPM_q_ivl_38712,
      c => LPM_d0_ivl_38729,
      clk => clk,
      r => LPM_q_ivl_38719
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3222
  SboxInst_U331: not_masked
    port map (
      a => LPM_q_ivl_6494,
      b => LPM_d0_ivl_6496
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4752
  SboxInst_U332: nor_HPC2
    port map (
      a => LPM_q_ivl_38675,
      b => LPM_q_ivl_38682,
      c => LPM_d0_ivl_38699,
      clk => clk,
      r => LPM_q_ivl_38689
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3221
  SboxInst_U333: not_masked
    port map (
      a => LPM_q_ivl_6487,
      b => LPM_d0_ivl_6489
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4751
  SboxInst_U334: nor_HPC2
    port map (
      a => LPM_q_ivl_38645,
      b => LPM_q_ivl_38652,
      c => LPM_d0_ivl_38669,
      clk => clk,
      r => LPM_q_ivl_38659
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3220
  SboxInst_U335: not_masked
    port map (
      a => LPM_q_ivl_6480,
      b => LPM_d0_ivl_6482
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4750
  SboxInst_U336: nor_HPC2
    port map (
      a => LPM_q_ivl_38615,
      b => LPM_q_ivl_38622,
      c => LPM_d0_ivl_38639,
      clk => clk,
      r => LPM_q_ivl_38629
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3219
  SboxInst_U337: not_masked
    port map (
      a => LPM_q_ivl_6473,
      b => LPM_d0_ivl_6475
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4749
  SboxInst_U338: nor_HPC2
    port map (
      a => LPM_q_ivl_38585,
      b => LPM_q_ivl_38592,
      c => LPM_d0_ivl_38609,
      clk => clk,
      r => LPM_q_ivl_38599
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3218
  SboxInst_U339: not_masked
    port map (
      a => LPM_q_ivl_6466,
      b => LPM_d0_ivl_6468
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4933
  SboxInst_U34: and_HPC2
    port map (
      a => LPM_q_ivl_43979,
      b => LPM_q_ivl_43988,
      c => LPM_d0_ivl_44005,
      clk => clk,
      r => LPM_q_ivl_43995
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4748
  SboxInst_U340: nor_HPC2
    port map (
      a => LPM_q_ivl_38555,
      b => LPM_q_ivl_38562,
      c => LPM_d0_ivl_38579,
      clk => clk,
      r => LPM_q_ivl_38569
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3217
  SboxInst_U341: not_masked
    port map (
      a => LPM_q_ivl_6459,
      b => LPM_d0_ivl_6461
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4747
  SboxInst_U342: nor_HPC2
    port map (
      a => LPM_q_ivl_38525,
      b => LPM_q_ivl_38532,
      c => LPM_d0_ivl_38549,
      clk => clk,
      r => LPM_q_ivl_38539
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3216
  SboxInst_U343: not_masked
    port map (
      a => LPM_q_ivl_6452,
      b => LPM_d0_ivl_6454
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4746
  SboxInst_U344: nor_HPC2
    port map (
      a => LPM_q_ivl_38495,
      b => LPM_q_ivl_38502,
      c => LPM_d0_ivl_38519,
      clk => clk,
      r => LPM_q_ivl_38509
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3215
  SboxInst_U345: not_masked
    port map (
      a => LPM_q_ivl_6445,
      b => LPM_d0_ivl_6447
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4745
  SboxInst_U346: nor_HPC2
    port map (
      a => LPM_q_ivl_38465,
      b => LPM_q_ivl_38472,
      c => LPM_d0_ivl_38489,
      clk => clk,
      r => LPM_q_ivl_38479
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3214
  SboxInst_U347: not_masked
    port map (
      a => LPM_q_ivl_6438,
      b => LPM_d0_ivl_6440
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4744
  SboxInst_U348: nor_HPC2
    port map (
      a => LPM_q_ivl_38435,
      b => LPM_q_ivl_38442,
      c => LPM_d0_ivl_38459,
      clk => clk,
      r => LPM_q_ivl_38449
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3213
  SboxInst_U349: not_masked
    port map (
      a => LPM_q_ivl_6431,
      b => LPM_d0_ivl_6433
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3338
  SboxInst_U35: not_masked
    port map (
      a => LPM_q_ivl_7528,
      b => LPM_d0_ivl_7530
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4743
  SboxInst_U350: nor_HPC2
    port map (
      a => LPM_q_ivl_38405,
      b => LPM_q_ivl_38412,
      c => LPM_d0_ivl_38429,
      clk => clk,
      r => LPM_q_ivl_38419
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3212
  SboxInst_U351: not_masked
    port map (
      a => LPM_q_ivl_6424,
      b => LPM_d0_ivl_6426
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4742
  SboxInst_U352: nor_HPC2
    port map (
      a => LPM_q_ivl_38375,
      b => LPM_q_ivl_38382,
      c => LPM_d0_ivl_38399,
      clk => clk,
      r => LPM_q_ivl_38389
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3211
  SboxInst_U353: not_masked
    port map (
      a => LPM_q_ivl_6417,
      b => LPM_d0_ivl_6419
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4741
  SboxInst_U354: nor_HPC2
    port map (
      a => LPM_q_ivl_38345,
      b => LPM_q_ivl_38352,
      c => LPM_d0_ivl_38369,
      clk => clk,
      r => LPM_q_ivl_38359
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3210
  SboxInst_U355: not_masked
    port map (
      a => LPM_q_ivl_6410,
      b => LPM_d0_ivl_6412
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4740
  SboxInst_U356: nor_HPC2
    port map (
      a => LPM_q_ivl_38315,
      b => LPM_q_ivl_38322,
      c => LPM_d0_ivl_38339,
      clk => clk,
      r => LPM_q_ivl_38329
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3209
  SboxInst_U357: not_masked
    port map (
      a => LPM_q_ivl_6403,
      b => LPM_d0_ivl_6405
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4739
  SboxInst_U358: nor_HPC2
    port map (
      a => LPM_q_ivl_38285,
      b => LPM_q_ivl_38292,
      c => LPM_d0_ivl_38309,
      clk => clk,
      r => LPM_q_ivl_38299
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3208
  SboxInst_U359: not_masked
    port map (
      a => LPM_q_ivl_6396,
      b => LPM_d0_ivl_6398
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4932
  SboxInst_U36: and_HPC2
    port map (
      a => LPM_q_ivl_43949,
      b => LPM_q_ivl_43958,
      c => LPM_d0_ivl_43975,
      clk => clk,
      r => LPM_q_ivl_43965
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4738
  SboxInst_U360: nor_HPC2
    port map (
      a => LPM_q_ivl_38255,
      b => LPM_q_ivl_38262,
      c => LPM_d0_ivl_38279,
      clk => clk,
      r => LPM_q_ivl_38269
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3207
  SboxInst_U361: not_masked
    port map (
      a => LPM_q_ivl_6389,
      b => LPM_d0_ivl_6391
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4737
  SboxInst_U362: nor_HPC2
    port map (
      a => LPM_q_ivl_38225,
      b => LPM_q_ivl_38232,
      c => LPM_d0_ivl_38249,
      clk => clk,
      r => LPM_q_ivl_38239
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3206
  SboxInst_U363: not_masked
    port map (
      a => LPM_q_ivl_6382,
      b => LPM_d0_ivl_6384
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4736
  SboxInst_U364: nor_HPC2
    port map (
      a => LPM_q_ivl_38195,
      b => LPM_q_ivl_38202,
      c => LPM_d0_ivl_38219,
      clk => clk,
      r => LPM_q_ivl_38209
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3205
  SboxInst_U365: not_masked
    port map (
      a => LPM_q_ivl_6375,
      b => LPM_d0_ivl_6377
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4735
  SboxInst_U366: nor_HPC2
    port map (
      a => LPM_q_ivl_38165,
      b => LPM_q_ivl_38172,
      c => LPM_d0_ivl_38189,
      clk => clk,
      r => LPM_q_ivl_38179
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3204
  SboxInst_U367: not_masked
    port map (
      a => LPM_q_ivl_6368,
      b => LPM_d0_ivl_6370
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4734
  SboxInst_U368: nor_HPC2
    port map (
      a => LPM_q_ivl_38135,
      b => LPM_q_ivl_38142,
      c => LPM_d0_ivl_38159,
      clk => clk,
      r => LPM_q_ivl_38149
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3203
  SboxInst_U369: not_masked
    port map (
      a => LPM_q_ivl_6361,
      b => LPM_d0_ivl_6363
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3337
  SboxInst_U37: not_masked
    port map (
      a => LPM_q_ivl_7519,
      b => LPM_d0_ivl_7521
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4733
  SboxInst_U370: nor_HPC2
    port map (
      a => LPM_q_ivl_38105,
      b => LPM_q_ivl_38112,
      c => LPM_d0_ivl_38129,
      clk => clk,
      r => LPM_q_ivl_38119
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3202
  SboxInst_U371: not_masked
    port map (
      a => LPM_q_ivl_6354,
      b => LPM_d0_ivl_6356
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4732
  SboxInst_U372: nor_HPC2
    port map (
      a => LPM_q_ivl_38075,
      b => LPM_q_ivl_38082,
      c => LPM_d0_ivl_38099,
      clk => clk,
      r => LPM_q_ivl_38089
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3201
  SboxInst_U373: not_masked
    port map (
      a => LPM_q_ivl_6347,
      b => LPM_d0_ivl_6349
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4731
  SboxInst_U374: nor_HPC2
    port map (
      a => LPM_q_ivl_38045,
      b => LPM_q_ivl_38052,
      c => LPM_d0_ivl_38069,
      clk => clk,
      r => LPM_q_ivl_38059
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3200
  SboxInst_U375: not_masked
    port map (
      a => LPM_q_ivl_6340,
      b => LPM_d0_ivl_6342
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4730
  SboxInst_U376: nor_HPC2
    port map (
      a => LPM_q_ivl_38015,
      b => LPM_q_ivl_38022,
      c => LPM_d0_ivl_38039,
      clk => clk,
      r => LPM_q_ivl_38029
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3199
  SboxInst_U377: not_masked
    port map (
      a => LPM_q_ivl_6333,
      b => LPM_d0_ivl_6335
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4729
  SboxInst_U378: nor_HPC2
    port map (
      a => LPM_q_ivl_37985,
      b => LPM_q_ivl_37992,
      c => LPM_d0_ivl_38009,
      clk => clk,
      r => LPM_q_ivl_37999
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3198
  SboxInst_U379: not_masked
    port map (
      a => LPM_q_ivl_6326,
      b => LPM_d0_ivl_6328
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4931
  SboxInst_U38: and_HPC2
    port map (
      a => LPM_q_ivl_43919,
      b => LPM_q_ivl_43928,
      c => LPM_d0_ivl_43945,
      clk => clk,
      r => LPM_q_ivl_43935
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4728
  SboxInst_U380: nor_HPC2
    port map (
      a => LPM_q_ivl_37955,
      b => LPM_q_ivl_37962,
      c => LPM_d0_ivl_37979,
      clk => clk,
      r => LPM_q_ivl_37969
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3197
  SboxInst_U381: not_masked
    port map (
      a => LPM_q_ivl_6319,
      b => LPM_d0_ivl_6321
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4727
  SboxInst_U382: nor_HPC2
    port map (
      a => LPM_q_ivl_37925,
      b => LPM_q_ivl_37932,
      c => LPM_d0_ivl_37949,
      clk => clk,
      r => LPM_q_ivl_37939
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3196
  SboxInst_U383: not_masked
    port map (
      a => LPM_q_ivl_6312,
      b => LPM_d0_ivl_6314
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4726
  SboxInst_U384: nor_HPC2
    port map (
      a => LPM_q_ivl_37895,
      b => LPM_q_ivl_37902,
      c => LPM_d0_ivl_37919,
      clk => clk,
      r => LPM_q_ivl_37909
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3195
  SboxInst_U385: not_masked
    port map (
      a => LPM_q_ivl_6305,
      b => LPM_d0_ivl_6307
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4725
  SboxInst_U386: nor_HPC2
    port map (
      a => LPM_q_ivl_37865,
      b => LPM_q_ivl_37872,
      c => LPM_d0_ivl_37889,
      clk => clk,
      r => LPM_q_ivl_37879
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3194
  SboxInst_U387: not_masked
    port map (
      a => LPM_q_ivl_6298,
      b => LPM_d0_ivl_6300
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4724
  SboxInst_U388: nor_HPC2
    port map (
      a => LPM_q_ivl_37835,
      b => LPM_q_ivl_37842,
      c => LPM_d0_ivl_37859,
      clk => clk,
      r => LPM_q_ivl_37849
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3193
  SboxInst_U389: not_masked
    port map (
      a => LPM_q_ivl_6291,
      b => LPM_d0_ivl_6293
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3336
  SboxInst_U39: not_masked
    port map (
      a => LPM_q_ivl_7510,
      b => LPM_d0_ivl_7512
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4723
  SboxInst_U390: nor_HPC2
    port map (
      a => LPM_q_ivl_37805,
      b => LPM_q_ivl_37812,
      c => LPM_d0_ivl_37829,
      clk => clk,
      r => LPM_q_ivl_37819
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3192
  SboxInst_U391: not_masked
    port map (
      a => LPM_q_ivl_6284,
      b => LPM_d0_ivl_6286
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4722
  SboxInst_U392: nor_HPC2
    port map (
      a => LPM_q_ivl_37775,
      b => LPM_q_ivl_37782,
      c => LPM_d0_ivl_37799,
      clk => clk,
      r => LPM_q_ivl_37789
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3191
  SboxInst_U393: not_masked
    port map (
      a => LPM_q_ivl_6277,
      b => LPM_d0_ivl_6279
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4721
  SboxInst_U394: nor_HPC2
    port map (
      a => LPM_q_ivl_37745,
      b => LPM_q_ivl_37752,
      c => LPM_d0_ivl_37769,
      clk => clk,
      r => LPM_q_ivl_37759
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3190
  SboxInst_U395: not_masked
    port map (
      a => LPM_q_ivl_6270,
      b => LPM_d0_ivl_6272
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4720
  SboxInst_U396: nor_HPC2
    port map (
      a => LPM_q_ivl_37715,
      b => LPM_q_ivl_37722,
      c => LPM_d0_ivl_37739,
      clk => clk,
      r => LPM_q_ivl_37729
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3189
  SboxInst_U397: not_masked
    port map (
      a => LPM_q_ivl_6263,
      b => LPM_d0_ivl_6265
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4719
  SboxInst_U398: nor_HPC2
    port map (
      a => LPM_q_ivl_37685,
      b => LPM_q_ivl_37692,
      c => LPM_d0_ivl_37709,
      clk => clk,
      r => LPM_q_ivl_37699
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3188
  SboxInst_U399: not_masked
    port map (
      a => LPM_q_ivl_6256,
      b => LPM_d0_ivl_6258
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4948
  SboxInst_U4: and_HPC2
    port map (
      a => LPM_q_ivl_44429,
      b => LPM_q_ivl_44438,
      c => LPM_d0_ivl_44455,
      clk => clk,
      r => LPM_q_ivl_44445
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4930
  SboxInst_U40: and_HPC2
    port map (
      a => LPM_q_ivl_43889,
      b => LPM_q_ivl_43898,
      c => LPM_d0_ivl_43915,
      clk => clk,
      r => LPM_q_ivl_43905
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4718
  SboxInst_U400: nor_HPC2
    port map (
      a => LPM_q_ivl_37655,
      b => LPM_q_ivl_37662,
      c => LPM_d0_ivl_37679,
      clk => clk,
      r => LPM_q_ivl_37669
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3187
  SboxInst_U401: not_masked
    port map (
      a => LPM_q_ivl_6249,
      b => LPM_d0_ivl_6251
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4717
  SboxInst_U402: nor_HPC2
    port map (
      a => LPM_q_ivl_37625,
      b => LPM_q_ivl_37632,
      c => LPM_d0_ivl_37649,
      clk => clk,
      r => LPM_q_ivl_37639
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3186
  SboxInst_U403: not_masked
    port map (
      a => LPM_q_ivl_6242,
      b => LPM_d0_ivl_6244
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4716
  SboxInst_U404: nor_HPC2
    port map (
      a => LPM_q_ivl_37595,
      b => LPM_q_ivl_37602,
      c => LPM_d0_ivl_37619,
      clk => clk,
      r => LPM_q_ivl_37609
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3185
  SboxInst_U405: not_masked
    port map (
      a => LPM_q_ivl_6235,
      b => LPM_d0_ivl_6237
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4715
  SboxInst_U406: nor_HPC2
    port map (
      a => LPM_q_ivl_37565,
      b => LPM_q_ivl_37572,
      c => LPM_d0_ivl_37589,
      clk => clk,
      r => LPM_q_ivl_37579
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3184
  SboxInst_U407: not_masked
    port map (
      a => LPM_q_ivl_6228,
      b => LPM_d0_ivl_6230
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4714
  SboxInst_U408: nor_HPC2
    port map (
      a => LPM_q_ivl_37535,
      b => LPM_q_ivl_37542,
      c => LPM_d0_ivl_37559,
      clk => clk,
      r => LPM_q_ivl_37549
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3183
  SboxInst_U409: not_masked
    port map (
      a => LPM_q_ivl_6221,
      b => LPM_d0_ivl_6223
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3335
  SboxInst_U41: not_masked
    port map (
      a => LPM_q_ivl_7501,
      b => LPM_d0_ivl_7503
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4713
  SboxInst_U410: nor_HPC2
    port map (
      a => LPM_q_ivl_37505,
      b => LPM_q_ivl_37512,
      c => LPM_d0_ivl_37529,
      clk => clk,
      r => LPM_q_ivl_37519
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3182
  SboxInst_U411: not_masked
    port map (
      a => LPM_q_ivl_6214,
      b => LPM_d0_ivl_6216
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4712
  SboxInst_U412: nor_HPC2
    port map (
      a => LPM_q_ivl_37475,
      b => LPM_q_ivl_37482,
      c => LPM_d0_ivl_37499,
      clk => clk,
      r => LPM_q_ivl_37489
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3181
  SboxInst_U413: not_masked
    port map (
      a => LPM_q_ivl_6207,
      b => LPM_d0_ivl_6209
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4711
  SboxInst_U414: nor_HPC2
    port map (
      a => LPM_q_ivl_37445,
      b => LPM_q_ivl_37452,
      c => LPM_d0_ivl_37469,
      clk => clk,
      r => LPM_q_ivl_37459
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3180
  SboxInst_U415: not_masked
    port map (
      a => LPM_q_ivl_6200,
      b => LPM_d0_ivl_6202
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4710
  SboxInst_U416: nor_HPC2
    port map (
      a => LPM_q_ivl_37415,
      b => LPM_q_ivl_37422,
      c => LPM_d0_ivl_37439,
      clk => clk,
      r => LPM_q_ivl_37429
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3179
  SboxInst_U417: not_masked
    port map (
      a => LPM_q_ivl_6193,
      b => LPM_d0_ivl_6195
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4709
  SboxInst_U418: nor_HPC2
    port map (
      a => LPM_q_ivl_37385,
      b => LPM_q_ivl_37392,
      c => LPM_d0_ivl_37409,
      clk => clk,
      r => LPM_q_ivl_37399
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3178
  SboxInst_U419: not_masked
    port map (
      a => LPM_q_ivl_6186,
      b => LPM_d0_ivl_6188
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4929
  SboxInst_U42: and_HPC2
    port map (
      a => LPM_q_ivl_43859,
      b => LPM_q_ivl_43868,
      c => LPM_d0_ivl_43885,
      clk => clk,
      r => LPM_q_ivl_43875
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4708
  SboxInst_U420: nor_HPC2
    port map (
      a => LPM_q_ivl_37355,
      b => LPM_q_ivl_37362,
      c => LPM_d0_ivl_37379,
      clk => clk,
      r => LPM_q_ivl_37369
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3177
  SboxInst_U421: not_masked
    port map (
      a => LPM_q_ivl_6179,
      b => LPM_d0_ivl_6181
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4707
  SboxInst_U422: nor_HPC2
    port map (
      a => LPM_q_ivl_37325,
      b => LPM_q_ivl_37332,
      c => LPM_d0_ivl_37349,
      clk => clk,
      r => LPM_q_ivl_37339
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3176
  SboxInst_U423: not_masked
    port map (
      a => LPM_q_ivl_6172,
      b => LPM_d0_ivl_6174
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4706
  SboxInst_U424: nor_HPC2
    port map (
      a => LPM_q_ivl_37295,
      b => LPM_q_ivl_37302,
      c => LPM_d0_ivl_37319,
      clk => clk,
      r => LPM_q_ivl_37309
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3175
  SboxInst_U425: not_masked
    port map (
      a => LPM_q_ivl_6165,
      b => LPM_d0_ivl_6167
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4705
  SboxInst_U426: nor_HPC2
    port map (
      a => LPM_q_ivl_37265,
      b => LPM_q_ivl_37272,
      c => LPM_d0_ivl_37289,
      clk => clk,
      r => LPM_q_ivl_37279
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3174
  SboxInst_U427: not_masked
    port map (
      a => LPM_q_ivl_6158,
      b => LPM_d0_ivl_6160
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4704
  SboxInst_U428: nor_HPC2
    port map (
      a => LPM_q_ivl_37235,
      b => LPM_q_ivl_37242,
      c => LPM_d0_ivl_37259,
      clk => clk,
      r => LPM_q_ivl_37249
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3173
  SboxInst_U429: not_masked
    port map (
      a => LPM_q_ivl_6151,
      b => LPM_d0_ivl_6153
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3334
  SboxInst_U43: not_masked
    port map (
      a => LPM_q_ivl_7492,
      b => LPM_d0_ivl_7494
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4703
  SboxInst_U430: nor_HPC2
    port map (
      a => LPM_q_ivl_37205,
      b => LPM_q_ivl_37212,
      c => LPM_d0_ivl_37229,
      clk => clk,
      r => LPM_q_ivl_37219
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3172
  SboxInst_U431: not_masked
    port map (
      a => LPM_q_ivl_6144,
      b => LPM_d0_ivl_6146
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4702
  SboxInst_U432: nor_HPC2
    port map (
      a => LPM_q_ivl_37175,
      b => LPM_q_ivl_37182,
      c => LPM_d0_ivl_37199,
      clk => clk,
      r => LPM_q_ivl_37189
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3171
  SboxInst_U433: not_masked
    port map (
      a => LPM_q_ivl_6137,
      b => LPM_d0_ivl_6139
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4701
  SboxInst_U434: nor_HPC2
    port map (
      a => LPM_q_ivl_37145,
      b => LPM_q_ivl_37152,
      c => LPM_d0_ivl_37169,
      clk => clk,
      r => LPM_q_ivl_37159
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3170
  SboxInst_U435: not_masked
    port map (
      a => LPM_q_ivl_6130,
      b => LPM_d0_ivl_6132
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4700
  SboxInst_U436: nor_HPC2
    port map (
      a => LPM_q_ivl_37115,
      b => LPM_q_ivl_37122,
      c => LPM_d0_ivl_37139,
      clk => clk,
      r => LPM_q_ivl_37129
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3169
  SboxInst_U437: not_masked
    port map (
      a => LPM_q_ivl_6123,
      b => LPM_d0_ivl_6125
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4699
  SboxInst_U438: nor_HPC2
    port map (
      a => LPM_q_ivl_37085,
      b => LPM_q_ivl_37092,
      c => LPM_d0_ivl_37109,
      clk => clk,
      r => LPM_q_ivl_37099
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3168
  SboxInst_U439: not_masked
    port map (
      a => LPM_q_ivl_6116,
      b => LPM_d0_ivl_6118
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4928
  SboxInst_U44: and_HPC2
    port map (
      a => LPM_q_ivl_43829,
      b => LPM_q_ivl_43838,
      c => LPM_d0_ivl_43855,
      clk => clk,
      r => LPM_q_ivl_43845
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4698
  SboxInst_U440: nor_HPC2
    port map (
      a => LPM_q_ivl_37055,
      b => LPM_q_ivl_37062,
      c => LPM_d0_ivl_37079,
      clk => clk,
      r => LPM_q_ivl_37069
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3167
  SboxInst_U441: not_masked
    port map (
      a => LPM_q_ivl_6109,
      b => LPM_d0_ivl_6111
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4697
  SboxInst_U442: nor_HPC2
    port map (
      a => LPM_q_ivl_37025,
      b => LPM_q_ivl_37032,
      c => LPM_d0_ivl_37049,
      clk => clk,
      r => LPM_q_ivl_37039
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3166
  SboxInst_U443: not_masked
    port map (
      a => LPM_q_ivl_6102,
      b => LPM_d0_ivl_6104
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4696
  SboxInst_U444: nor_HPC2
    port map (
      a => LPM_q_ivl_36995,
      b => LPM_q_ivl_37002,
      c => LPM_d0_ivl_37019,
      clk => clk,
      r => LPM_q_ivl_37009
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3165
  SboxInst_U445: not_masked
    port map (
      a => LPM_q_ivl_6095,
      b => LPM_d0_ivl_6097
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4695
  SboxInst_U446: nor_HPC2
    port map (
      a => LPM_q_ivl_36965,
      b => LPM_q_ivl_36972,
      c => LPM_d0_ivl_36989,
      clk => clk,
      r => LPM_q_ivl_36979
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3164
  SboxInst_U447: not_masked
    port map (
      a => LPM_q_ivl_6088,
      b => LPM_d0_ivl_6090
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4694
  SboxInst_U448: nor_HPC2
    port map (
      a => LPM_q_ivl_36935,
      b => LPM_q_ivl_36942,
      c => LPM_d0_ivl_36959,
      clk => clk,
      r => LPM_q_ivl_36949
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4693
  SboxInst_U449: nor_HPC2
    port map (
      a => LPM_q_ivl_36905,
      b => LPM_q_ivl_36912,
      c => LPM_d0_ivl_36929,
      clk => clk,
      r => LPM_q_ivl_36919
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3333
  SboxInst_U45: not_masked
    port map (
      a => LPM_q_ivl_7483,
      b => LPM_d0_ivl_7485
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4692
  SboxInst_U450: nor_HPC2
    port map (
      a => LPM_q_ivl_36877,
      b => LPM_q_ivl_36884,
      c => LPM_d0_ivl_36901,
      clk => clk,
      r => LPM_q_ivl_36891
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4691
  SboxInst_U451: nor_HPC2
    port map (
      a => LPM_q_ivl_36849,
      b => LPM_q_ivl_36856,
      c => LPM_d0_ivl_36873,
      clk => clk,
      r => LPM_q_ivl_36863
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4690
  SboxInst_U452: nor_HPC2
    port map (
      a => LPM_q_ivl_36821,
      b => LPM_q_ivl_36828,
      c => LPM_d0_ivl_36845,
      clk => clk,
      r => LPM_q_ivl_36835
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4689
  SboxInst_U453: nor_HPC2
    port map (
      a => LPM_q_ivl_36793,
      b => LPM_q_ivl_36800,
      c => LPM_d0_ivl_36817,
      clk => clk,
      r => LPM_q_ivl_36807
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4688
  SboxInst_U454: nor_HPC2
    port map (
      a => LPM_q_ivl_36765,
      b => LPM_q_ivl_36772,
      c => LPM_d0_ivl_36789,
      clk => clk,
      r => LPM_q_ivl_36779
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4687
  SboxInst_U455: nor_HPC2
    port map (
      a => LPM_q_ivl_36737,
      b => LPM_q_ivl_36744,
      c => LPM_d0_ivl_36761,
      clk => clk,
      r => LPM_q_ivl_36751
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4686
  SboxInst_U456: nor_HPC2
    port map (
      a => LPM_q_ivl_36709,
      b => LPM_q_ivl_36716,
      c => LPM_d0_ivl_36733,
      clk => clk,
      r => LPM_q_ivl_36723
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4685
  SboxInst_U457: nor_HPC2
    port map (
      a => LPM_q_ivl_36681,
      b => LPM_q_ivl_36688,
      c => LPM_d0_ivl_36705,
      clk => clk,
      r => LPM_q_ivl_36695
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4684
  SboxInst_U458: nor_HPC2
    port map (
      a => LPM_q_ivl_36653,
      b => LPM_q_ivl_36660,
      c => LPM_d0_ivl_36677,
      clk => clk,
      r => LPM_q_ivl_36667
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4683
  SboxInst_U459: nor_HPC2
    port map (
      a => LPM_q_ivl_36625,
      b => LPM_q_ivl_36632,
      c => LPM_d0_ivl_36649,
      clk => clk,
      r => LPM_q_ivl_36639
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4927
  SboxInst_U46: and_HPC2
    port map (
      a => LPM_q_ivl_43799,
      b => LPM_q_ivl_43808,
      c => LPM_d0_ivl_43825,
      clk => clk,
      r => LPM_q_ivl_43815
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4682
  SboxInst_U460: nor_HPC2
    port map (
      a => LPM_q_ivl_36597,
      b => LPM_q_ivl_36604,
      c => LPM_d0_ivl_36621,
      clk => clk,
      r => LPM_q_ivl_36611
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4681
  SboxInst_U461: nor_HPC2
    port map (
      a => LPM_q_ivl_36569,
      b => LPM_q_ivl_36576,
      c => LPM_d0_ivl_36593,
      clk => clk,
      r => LPM_q_ivl_36583
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4680
  SboxInst_U462: nor_HPC2
    port map (
      a => LPM_q_ivl_36541,
      b => LPM_q_ivl_36548,
      c => LPM_d0_ivl_36565,
      clk => clk,
      r => LPM_q_ivl_36555
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4679
  SboxInst_U463: nor_HPC2
    port map (
      a => LPM_q_ivl_36513,
      b => LPM_q_ivl_36520,
      c => LPM_d0_ivl_36537,
      clk => clk,
      r => LPM_q_ivl_36527
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4678
  SboxInst_U464: nor_HPC2
    port map (
      a => LPM_q_ivl_36485,
      b => LPM_q_ivl_36492,
      c => LPM_d0_ivl_36509,
      clk => clk,
      r => LPM_q_ivl_36499
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4677
  SboxInst_U465: nor_HPC2
    port map (
      a => LPM_q_ivl_36457,
      b => LPM_q_ivl_36464,
      c => LPM_d0_ivl_36481,
      clk => clk,
      r => LPM_q_ivl_36471
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4676
  SboxInst_U466: nor_HPC2
    port map (
      a => LPM_q_ivl_36429,
      b => LPM_q_ivl_36436,
      c => LPM_d0_ivl_36453,
      clk => clk,
      r => LPM_q_ivl_36443
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4675
  SboxInst_U467: nor_HPC2
    port map (
      a => LPM_q_ivl_36401,
      b => LPM_q_ivl_36408,
      c => LPM_d0_ivl_36425,
      clk => clk,
      r => LPM_q_ivl_36415
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4674
  SboxInst_U468: nor_HPC2
    port map (
      a => LPM_q_ivl_36373,
      b => LPM_q_ivl_36380,
      c => LPM_d0_ivl_36397,
      clk => clk,
      r => LPM_q_ivl_36387
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4673
  SboxInst_U469: nor_HPC2
    port map (
      a => LPM_q_ivl_36345,
      b => LPM_q_ivl_36352,
      c => LPM_d0_ivl_36369,
      clk => clk,
      r => LPM_q_ivl_36359
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3332
  SboxInst_U47: not_masked
    port map (
      a => LPM_q_ivl_7474,
      b => LPM_d0_ivl_7476
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4672
  SboxInst_U470: nor_HPC2
    port map (
      a => LPM_q_ivl_36317,
      b => LPM_q_ivl_36324,
      c => LPM_d0_ivl_36341,
      clk => clk,
      r => LPM_q_ivl_36331
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4671
  SboxInst_U471: nor_HPC2
    port map (
      a => LPM_q_ivl_36289,
      b => LPM_q_ivl_36296,
      c => LPM_d0_ivl_36313,
      clk => clk,
      r => LPM_q_ivl_36303
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4670
  SboxInst_U472: nor_HPC2
    port map (
      a => LPM_q_ivl_36261,
      b => LPM_q_ivl_36268,
      c => LPM_d0_ivl_36285,
      clk => clk,
      r => LPM_q_ivl_36275
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4669
  SboxInst_U473: nor_HPC2
    port map (
      a => LPM_q_ivl_36233,
      b => LPM_q_ivl_36240,
      c => LPM_d0_ivl_36257,
      clk => clk,
      r => LPM_q_ivl_36247
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4668
  SboxInst_U474: nor_HPC2
    port map (
      a => LPM_q_ivl_36205,
      b => LPM_q_ivl_36212,
      c => LPM_d0_ivl_36229,
      clk => clk,
      r => LPM_q_ivl_36219
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4667
  SboxInst_U475: nor_HPC2
    port map (
      a => LPM_q_ivl_36177,
      b => LPM_q_ivl_36184,
      c => LPM_d0_ivl_36201,
      clk => clk,
      r => LPM_q_ivl_36191
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4666
  SboxInst_U476: nor_HPC2
    port map (
      a => LPM_q_ivl_36149,
      b => LPM_q_ivl_36156,
      c => LPM_d0_ivl_36173,
      clk => clk,
      r => LPM_q_ivl_36163
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4665
  SboxInst_U477: nor_HPC2
    port map (
      a => LPM_q_ivl_36121,
      b => LPM_q_ivl_36128,
      c => LPM_d0_ivl_36145,
      clk => clk,
      r => LPM_q_ivl_36135
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4664
  SboxInst_U478: nor_HPC2
    port map (
      a => LPM_q_ivl_36093,
      b => LPM_q_ivl_36100,
      c => LPM_d0_ivl_36117,
      clk => clk,
      r => LPM_q_ivl_36107
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4663
  SboxInst_U479: nor_HPC2
    port map (
      a => LPM_q_ivl_36065,
      b => LPM_q_ivl_36072,
      c => LPM_d0_ivl_36089,
      clk => clk,
      r => LPM_q_ivl_36079
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4926
  SboxInst_U48: and_HPC2
    port map (
      a => LPM_q_ivl_43769,
      b => LPM_q_ivl_43778,
      c => LPM_d0_ivl_43795,
      clk => clk,
      r => LPM_q_ivl_43785
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4662
  SboxInst_U480: nor_HPC2
    port map (
      a => LPM_q_ivl_36037,
      b => LPM_q_ivl_36044,
      c => LPM_d0_ivl_36061,
      clk => clk,
      r => LPM_q_ivl_36051
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4661
  SboxInst_U481: nor_HPC2
    port map (
      a => LPM_q_ivl_36009,
      b => LPM_q_ivl_36016,
      c => LPM_d0_ivl_36033,
      clk => clk,
      r => LPM_q_ivl_36023
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4660
  SboxInst_U482: nor_HPC2
    port map (
      a => LPM_q_ivl_35981,
      b => LPM_q_ivl_35988,
      c => LPM_d0_ivl_36005,
      clk => clk,
      r => LPM_q_ivl_35995
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4659
  SboxInst_U483: nor_HPC2
    port map (
      a => LPM_q_ivl_35953,
      b => LPM_q_ivl_35960,
      c => LPM_d0_ivl_35977,
      clk => clk,
      r => LPM_q_ivl_35967
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4658
  SboxInst_U484: nor_HPC2
    port map (
      a => LPM_q_ivl_35925,
      b => LPM_q_ivl_35932,
      c => LPM_d0_ivl_35949,
      clk => clk,
      r => LPM_q_ivl_35939
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4657
  SboxInst_U485: nor_HPC2
    port map (
      a => LPM_q_ivl_35897,
      b => LPM_q_ivl_35904,
      c => LPM_d0_ivl_35921,
      clk => clk,
      r => LPM_q_ivl_35911
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4656
  SboxInst_U486: nor_HPC2
    port map (
      a => LPM_q_ivl_35869,
      b => LPM_q_ivl_35876,
      c => LPM_d0_ivl_35893,
      clk => clk,
      r => LPM_q_ivl_35883
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4655
  SboxInst_U487: nor_HPC2
    port map (
      a => LPM_q_ivl_35841,
      b => LPM_q_ivl_35848,
      c => LPM_d0_ivl_35865,
      clk => clk,
      r => LPM_q_ivl_35855
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4654
  SboxInst_U488: nor_HPC2
    port map (
      a => LPM_q_ivl_35813,
      b => LPM_q_ivl_35820,
      c => LPM_d0_ivl_35837,
      clk => clk,
      r => LPM_q_ivl_35827
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4653
  SboxInst_U489: nor_HPC2
    port map (
      a => LPM_q_ivl_35785,
      b => LPM_q_ivl_35792,
      c => LPM_d0_ivl_35809,
      clk => clk,
      r => LPM_q_ivl_35799
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3331
  SboxInst_U49: not_masked
    port map (
      a => LPM_q_ivl_7465,
      b => LPM_d0_ivl_7467
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4652
  SboxInst_U490: nor_HPC2
    port map (
      a => LPM_q_ivl_35757,
      b => LPM_q_ivl_35764,
      c => LPM_d0_ivl_35781,
      clk => clk,
      r => LPM_q_ivl_35771
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4651
  SboxInst_U491: nor_HPC2
    port map (
      a => LPM_q_ivl_35729,
      b => LPM_q_ivl_35736,
      c => LPM_d0_ivl_35753,
      clk => clk,
      r => LPM_q_ivl_35743
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4650
  SboxInst_U492: nor_HPC2
    port map (
      a => LPM_q_ivl_35701,
      b => LPM_q_ivl_35708,
      c => LPM_d0_ivl_35725,
      clk => clk,
      r => LPM_q_ivl_35715
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4649
  SboxInst_U493: nor_HPC2
    port map (
      a => LPM_q_ivl_35673,
      b => LPM_q_ivl_35680,
      c => LPM_d0_ivl_35697,
      clk => clk,
      r => LPM_q_ivl_35687
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4648
  SboxInst_U494: nor_HPC2
    port map (
      a => LPM_q_ivl_35645,
      b => LPM_q_ivl_35652,
      c => LPM_d0_ivl_35669,
      clk => clk,
      r => LPM_q_ivl_35659
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4647
  SboxInst_U495: nor_HPC2
    port map (
      a => LPM_q_ivl_35617,
      b => LPM_q_ivl_35624,
      c => LPM_d0_ivl_35641,
      clk => clk,
      r => LPM_q_ivl_35631
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4646
  SboxInst_U496: nor_HPC2
    port map (
      a => LPM_q_ivl_35589,
      b => LPM_q_ivl_35596,
      c => LPM_d0_ivl_35613,
      clk => clk,
      r => LPM_q_ivl_35603
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4645
  SboxInst_U497: nor_HPC2
    port map (
      a => LPM_q_ivl_35561,
      b => LPM_q_ivl_35568,
      c => LPM_d0_ivl_35585,
      clk => clk,
      r => LPM_q_ivl_35575
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4644
  SboxInst_U498: nor_HPC2
    port map (
      a => LPM_q_ivl_35533,
      b => LPM_q_ivl_35540,
      c => LPM_d0_ivl_35557,
      clk => clk,
      r => LPM_q_ivl_35547
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4643
  SboxInst_U499: nor_HPC2
    port map (
      a => LPM_q_ivl_35505,
      b => LPM_q_ivl_35512,
      c => LPM_d0_ivl_35529,
      clk => clk,
      r => LPM_q_ivl_35519
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3353
  SboxInst_U5: not_masked
    port map (
      a => LPM_q_ivl_7663,
      b => LPM_d0_ivl_7665
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4925
  SboxInst_U50: and_HPC2
    port map (
      a => LPM_q_ivl_43739,
      b => LPM_q_ivl_43748,
      c => LPM_d0_ivl_43765,
      clk => clk,
      r => LPM_q_ivl_43755
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4642
  SboxInst_U500: nor_HPC2
    port map (
      a => LPM_q_ivl_35477,
      b => LPM_q_ivl_35484,
      c => LPM_d0_ivl_35501,
      clk => clk,
      r => LPM_q_ivl_35491
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4641
  SboxInst_U501: nor_HPC2
    port map (
      a => LPM_q_ivl_35449,
      b => LPM_q_ivl_35456,
      c => LPM_d0_ivl_35473,
      clk => clk,
      r => LPM_q_ivl_35463
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4640
  SboxInst_U502: nor_HPC2
    port map (
      a => LPM_q_ivl_35419,
      b => LPM_q_ivl_35426,
      c => LPM_d0_ivl_35443,
      clk => clk,
      r => LPM_q_ivl_35433
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4639
  SboxInst_U503: nor_HPC2
    port map (
      a => LPM_q_ivl_35391,
      b => LPM_q_ivl_35398,
      c => LPM_d0_ivl_35415,
      clk => clk,
      r => LPM_q_ivl_35405
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4638
  SboxInst_U504: nor_HPC2
    port map (
      a => LPM_q_ivl_35363,
      b => LPM_q_ivl_35370,
      c => LPM_d0_ivl_35387,
      clk => clk,
      r => LPM_q_ivl_35377
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4637
  SboxInst_U505: nor_HPC2
    port map (
      a => LPM_q_ivl_35335,
      b => LPM_q_ivl_35342,
      c => LPM_d0_ivl_35359,
      clk => clk,
      r => LPM_q_ivl_35349
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4636
  SboxInst_U506: nor_HPC2
    port map (
      a => LPM_q_ivl_35307,
      b => LPM_q_ivl_35314,
      c => LPM_d0_ivl_35331,
      clk => clk,
      r => LPM_q_ivl_35321
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4635
  SboxInst_U507: nor_HPC2
    port map (
      a => LPM_q_ivl_35279,
      b => LPM_q_ivl_35286,
      c => LPM_d0_ivl_35303,
      clk => clk,
      r => LPM_q_ivl_35293
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4634
  SboxInst_U508: nor_HPC2
    port map (
      a => LPM_q_ivl_35251,
      b => LPM_q_ivl_35258,
      c => LPM_d0_ivl_35275,
      clk => clk,
      r => LPM_q_ivl_35265
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4633
  SboxInst_U509: nor_HPC2
    port map (
      a => LPM_q_ivl_35223,
      b => LPM_q_ivl_35230,
      c => LPM_d0_ivl_35247,
      clk => clk,
      r => LPM_q_ivl_35237
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3330
  SboxInst_U51: not_masked
    port map (
      a => LPM_q_ivl_7456,
      b => LPM_d0_ivl_7458
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4632
  SboxInst_U510: nor_HPC2
    port map (
      a => LPM_q_ivl_35195,
      b => LPM_q_ivl_35202,
      c => LPM_d0_ivl_35219,
      clk => clk,
      r => LPM_q_ivl_35209
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4631
  SboxInst_U511: nor_HPC2
    port map (
      a => LPM_q_ivl_35167,
      b => LPM_q_ivl_35174,
      c => LPM_d0_ivl_35191,
      clk => clk,
      r => LPM_q_ivl_35181
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4630
  SboxInst_U512: nor_HPC2
    port map (
      a => LPM_q_ivl_35139,
      b => LPM_q_ivl_35146,
      c => LPM_d0_ivl_35163,
      clk => clk,
      r => LPM_q_ivl_35153
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4924
  SboxInst_U52: and_HPC2
    port map (
      a => LPM_q_ivl_43709,
      b => LPM_q_ivl_43718,
      c => LPM_d0_ivl_43735,
      clk => clk,
      r => LPM_q_ivl_43725
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3329
  SboxInst_U53: not_masked
    port map (
      a => LPM_q_ivl_7447,
      b => LPM_d0_ivl_7449
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4923
  SboxInst_U54: and_HPC2
    port map (
      a => LPM_q_ivl_43681,
      b => LPM_q_ivl_43688,
      c => LPM_d0_ivl_43705,
      clk => clk,
      r => LPM_q_ivl_43695
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3328
  SboxInst_U55: not_masked
    port map (
      a => LPM_q_ivl_7438,
      b => LPM_d0_ivl_7440
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4922
  SboxInst_U56: and_HPC2
    port map (
      a => LPM_q_ivl_43653,
      b => LPM_q_ivl_43660,
      c => LPM_d0_ivl_43677,
      clk => clk,
      r => LPM_q_ivl_43667
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3327
  SboxInst_U57: not_masked
    port map (
      a => LPM_q_ivl_7429,
      b => LPM_d0_ivl_7431
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4921
  SboxInst_U58: and_HPC2
    port map (
      a => LPM_q_ivl_43625,
      b => LPM_q_ivl_43632,
      c => LPM_d0_ivl_43649,
      clk => clk,
      r => LPM_q_ivl_43639
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3326
  SboxInst_U59: not_masked
    port map (
      a => LPM_q_ivl_7420,
      b => LPM_d0_ivl_7422
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4947
  SboxInst_U6: and_HPC2
    port map (
      a => LPM_q_ivl_44399,
      b => LPM_q_ivl_44408,
      c => LPM_d0_ivl_44425,
      clk => clk,
      r => LPM_q_ivl_44415
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4920
  SboxInst_U60: and_HPC2
    port map (
      a => LPM_q_ivl_43597,
      b => LPM_q_ivl_43604,
      c => LPM_d0_ivl_43621,
      clk => clk,
      r => LPM_q_ivl_43611
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3325
  SboxInst_U61: not_masked
    port map (
      a => LPM_q_ivl_7411,
      b => LPM_d0_ivl_7413
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4919
  SboxInst_U62: and_HPC2
    port map (
      a => LPM_q_ivl_43569,
      b => LPM_q_ivl_43576,
      c => LPM_d0_ivl_43593,
      clk => clk,
      r => LPM_q_ivl_43583
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3324
  SboxInst_U63: not_masked
    port map (
      a => LPM_q_ivl_7402,
      b => LPM_d0_ivl_7404
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4918
  SboxInst_U64: and_HPC2
    port map (
      a => LPM_q_ivl_43541,
      b => LPM_q_ivl_43548,
      c => LPM_d0_ivl_43565,
      clk => clk,
      r => LPM_q_ivl_43555
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3323
  SboxInst_U65: not_masked
    port map (
      a => LPM_q_ivl_7393,
      b => LPM_d0_ivl_7395
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4917
  SboxInst_U66: and_HPC2
    port map (
      a => LPM_q_ivl_43513,
      b => LPM_q_ivl_43520,
      c => LPM_d0_ivl_43537,
      clk => clk,
      r => LPM_q_ivl_43527
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3322
  SboxInst_U67: not_masked
    port map (
      a => LPM_q_ivl_7384,
      b => LPM_d0_ivl_7386
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4916
  SboxInst_U68: and_HPC2
    port map (
      a => LPM_q_ivl_43485,
      b => LPM_q_ivl_43492,
      c => LPM_d0_ivl_43509,
      clk => clk,
      r => LPM_q_ivl_43499
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3321
  SboxInst_U69: not_masked
    port map (
      a => LPM_q_ivl_7375,
      b => LPM_d0_ivl_7377
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3352
  SboxInst_U7: not_masked
    port map (
      a => LPM_q_ivl_7654,
      b => LPM_d0_ivl_7656
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4915
  SboxInst_U70: and_HPC2
    port map (
      a => LPM_q_ivl_43457,
      b => LPM_q_ivl_43464,
      c => LPM_d0_ivl_43481,
      clk => clk,
      r => LPM_q_ivl_43471
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3320
  SboxInst_U71: not_masked
    port map (
      a => LPM_q_ivl_7366,
      b => LPM_d0_ivl_7368
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4914
  SboxInst_U72: and_HPC2
    port map (
      a => LPM_q_ivl_43429,
      b => LPM_q_ivl_43436,
      c => LPM_d0_ivl_43453,
      clk => clk,
      r => LPM_q_ivl_43443
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3319
  SboxInst_U73: not_masked
    port map (
      a => LPM_q_ivl_7357,
      b => LPM_d0_ivl_7359
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4913
  SboxInst_U74: and_HPC2
    port map (
      a => LPM_q_ivl_43401,
      b => LPM_q_ivl_43408,
      c => LPM_d0_ivl_43425,
      clk => clk,
      r => LPM_q_ivl_43415
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3318
  SboxInst_U75: not_masked
    port map (
      a => LPM_q_ivl_7348,
      b => LPM_d0_ivl_7350
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4912
  SboxInst_U76: and_HPC2
    port map (
      a => LPM_q_ivl_43373,
      b => LPM_q_ivl_43380,
      c => LPM_d0_ivl_43397,
      clk => clk,
      r => LPM_q_ivl_43387
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3317
  SboxInst_U77: not_masked
    port map (
      a => LPM_q_ivl_7339,
      b => LPM_d0_ivl_7341
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4911
  SboxInst_U78: and_HPC2
    port map (
      a => LPM_q_ivl_43345,
      b => LPM_q_ivl_43352,
      c => LPM_d0_ivl_43369,
      clk => clk,
      r => LPM_q_ivl_43359
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3316
  SboxInst_U79: not_masked
    port map (
      a => LPM_q_ivl_7330,
      b => LPM_d0_ivl_7332
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4946
  SboxInst_U8: and_HPC2
    port map (
      a => LPM_q_ivl_44369,
      b => LPM_q_ivl_44378,
      c => LPM_d0_ivl_44395,
      clk => clk,
      r => LPM_q_ivl_44385
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4910
  SboxInst_U80: and_HPC2
    port map (
      a => LPM_q_ivl_43317,
      b => LPM_q_ivl_43324,
      c => LPM_d0_ivl_43341,
      clk => clk,
      r => LPM_q_ivl_43331
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3315
  SboxInst_U81: not_masked
    port map (
      a => LPM_q_ivl_7321,
      b => LPM_d0_ivl_7323
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4909
  SboxInst_U82: and_HPC2
    port map (
      a => LPM_q_ivl_43289,
      b => LPM_q_ivl_43296,
      c => LPM_d0_ivl_43313,
      clk => clk,
      r => LPM_q_ivl_43303
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3314
  SboxInst_U83: not_masked
    port map (
      a => LPM_q_ivl_7312,
      b => LPM_d0_ivl_7314
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4908
  SboxInst_U84: and_HPC2
    port map (
      a => LPM_q_ivl_43261,
      b => LPM_q_ivl_43268,
      c => LPM_d0_ivl_43285,
      clk => clk,
      r => LPM_q_ivl_43275
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3313
  SboxInst_U85: not_masked
    port map (
      a => LPM_q_ivl_7303,
      b => LPM_d0_ivl_7305
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4907
  SboxInst_U86: and_HPC2
    port map (
      a => LPM_q_ivl_43233,
      b => LPM_q_ivl_43240,
      c => LPM_d0_ivl_43257,
      clk => clk,
      r => LPM_q_ivl_43247
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3312
  SboxInst_U87: not_masked
    port map (
      a => LPM_q_ivl_7294,
      b => LPM_d0_ivl_7296
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4906
  SboxInst_U88: and_HPC2
    port map (
      a => LPM_q_ivl_43205,
      b => LPM_q_ivl_43212,
      c => LPM_d0_ivl_43229,
      clk => clk,
      r => LPM_q_ivl_43219
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3311
  SboxInst_U89: not_masked
    port map (
      a => LPM_q_ivl_7285,
      b => LPM_d0_ivl_7287
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3351
  SboxInst_U9: not_masked
    port map (
      a => LPM_q_ivl_7645,
      b => LPM_d0_ivl_7647
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4905
  SboxInst_U90: and_HPC2
    port map (
      a => LPM_q_ivl_43177,
      b => LPM_q_ivl_43184,
      c => LPM_d0_ivl_43201,
      clk => clk,
      r => LPM_q_ivl_43191
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3310
  SboxInst_U91: not_masked
    port map (
      a => LPM_q_ivl_7276,
      b => LPM_d0_ivl_7278
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4904
  SboxInst_U92: and_HPC2
    port map (
      a => LPM_q_ivl_43149,
      b => LPM_q_ivl_43156,
      c => LPM_d0_ivl_43173,
      clk => clk,
      r => LPM_q_ivl_43163
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3309
  SboxInst_U93: not_masked
    port map (
      a => LPM_q_ivl_7267,
      b => LPM_d0_ivl_7269
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4903
  SboxInst_U94: and_HPC2
    port map (
      a => LPM_q_ivl_43121,
      b => LPM_q_ivl_43128,
      c => LPM_d0_ivl_43145,
      clk => clk,
      r => LPM_q_ivl_43135
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3308
  SboxInst_U95: not_masked
    port map (
      a => LPM_q_ivl_7258,
      b => LPM_d0_ivl_7260
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4902
  SboxInst_U96: and_HPC2
    port map (
      a => LPM_q_ivl_43093,
      b => LPM_q_ivl_43100,
      c => LPM_d0_ivl_43117,
      clk => clk,
      r => LPM_q_ivl_43107
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3307
  SboxInst_U97: not_masked
    port map (
      a => LPM_q_ivl_7249,
      b => LPM_d0_ivl_7251
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4901
  SboxInst_U98: and_HPC2
    port map (
      a => LPM_q_ivl_43065,
      b => LPM_q_ivl_43072,
      c => LPM_d0_ivl_43089,
      clk => clk,
      r => LPM_q_ivl_43079
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3306
  SboxInst_U99: not_masked
    port map (
      a => LPM_q_ivl_7240,
      b => LPM_d0_ivl_7242
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2940
  U3097: xor_HPC2
    port map (
      a => LPM_q_ivl_7,
      b => LPM_q_ivl_18,
      c => LPM_d0_ivl_28
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2941
  U3098: xor_HPC2
    port map (
      a => LPM_q_ivl_36,
      b => LPM_q_ivl_47,
      c => LPM_d0_ivl_57
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2942
  U3099: xor_HPC2
    port map (
      a => LPM_q_ivl_65,
      b => LPM_q_ivl_76,
      c => LPM_d0_ivl_86
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2943
  U3100: xor_HPC2
    port map (
      a => LPM_q_ivl_94,
      b => LPM_q_ivl_105,
      c => LPM_d0_ivl_115
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2944
  U3101: xor_HPC2
    port map (
      a => LPM_q_ivl_123,
      b => LPM_q_ivl_134,
      c => LPM_d0_ivl_144
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2945
  U3102: xor_HPC2
    port map (
      a => LPM_q_ivl_152,
      b => LPM_q_ivl_163,
      c => LPM_d0_ivl_173
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2946
  U3103: xor_HPC2
    port map (
      a => LPM_q_ivl_181,
      b => LPM_q_ivl_192,
      c => LPM_d0_ivl_202
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2947
  U3104: xor_HPC2
    port map (
      a => LPM_q_ivl_210,
      b => LPM_q_ivl_221,
      c => LPM_d0_ivl_231
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2948
  U3105: xor_HPC2
    port map (
      a => LPM_q_ivl_239,
      b => LPM_q_ivl_250,
      c => LPM_d0_ivl_260
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2949
  U3106: xor_HPC2
    port map (
      a => LPM_q_ivl_268,
      b => LPM_q_ivl_279,
      c => LPM_d0_ivl_289
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2950
  U3107: xor_HPC2
    port map (
      a => LPM_q_ivl_297,
      b => LPM_q_ivl_308,
      c => LPM_d0_ivl_318
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2951
  U3108: xor_HPC2
    port map (
      a => LPM_q_ivl_326,
      b => LPM_q_ivl_337,
      c => LPM_d0_ivl_347
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2952
  U3109: xor_HPC2
    port map (
      a => LPM_q_ivl_355,
      b => LPM_q_ivl_366,
      c => LPM_d0_ivl_376
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2953
  U3110: xor_HPC2
    port map (
      a => LPM_q_ivl_384,
      b => LPM_q_ivl_395,
      c => LPM_d0_ivl_405
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2954
  U3111: xor_HPC2
    port map (
      a => LPM_q_ivl_413,
      b => LPM_q_ivl_424,
      c => LPM_d0_ivl_434
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2955
  U3112: xor_HPC2
    port map (
      a => LPM_q_ivl_442,
      b => LPM_q_ivl_453,
      c => LPM_d0_ivl_463
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2956
  U3113: xor_HPC2
    port map (
      a => LPM_q_ivl_471,
      b => LPM_q_ivl_482,
      c => LPM_d0_ivl_492
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2957
  U3114: xor_HPC2
    port map (
      a => LPM_q_ivl_500,
      b => LPM_q_ivl_511,
      c => LPM_d0_ivl_521
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2958
  U3115: xor_HPC2
    port map (
      a => LPM_q_ivl_529,
      b => LPM_q_ivl_540,
      c => LPM_d0_ivl_550
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2959
  U3116: xor_HPC2
    port map (
      a => LPM_q_ivl_558,
      b => LPM_q_ivl_569,
      c => LPM_d0_ivl_579
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2960
  U3117: xor_HPC2
    port map (
      a => LPM_q_ivl_587,
      b => LPM_q_ivl_598,
      c => LPM_d0_ivl_608
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2961
  U3118: xor_HPC2
    port map (
      a => LPM_q_ivl_616,
      b => LPM_q_ivl_627,
      c => LPM_d0_ivl_637
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2962
  U3119: xor_HPC2
    port map (
      a => LPM_q_ivl_645,
      b => LPM_q_ivl_656,
      c => LPM_d0_ivl_666
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2963
  U3120: xor_HPC2
    port map (
      a => LPM_q_ivl_674,
      b => LPM_q_ivl_685,
      c => LPM_d0_ivl_695
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2964
  U3121: xor_HPC2
    port map (
      a => LPM_q_ivl_703,
      b => LPM_q_ivl_714,
      c => LPM_d0_ivl_724
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2965
  U3122: xor_HPC2
    port map (
      a => LPM_q_ivl_732,
      b => LPM_q_ivl_743,
      c => LPM_d0_ivl_753
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2966
  U3123: xor_HPC2
    port map (
      a => LPM_q_ivl_761,
      b => LPM_q_ivl_772,
      c => LPM_d0_ivl_782
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2967
  U3124: xor_HPC2
    port map (
      a => LPM_q_ivl_790,
      b => LPM_q_ivl_801,
      c => LPM_d0_ivl_811
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2968
  U3125: xor_HPC2
    port map (
      a => LPM_q_ivl_819,
      b => LPM_q_ivl_830,
      c => LPM_d0_ivl_840
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2969
  U3126: xor_HPC2
    port map (
      a => LPM_q_ivl_848,
      b => LPM_q_ivl_859,
      c => LPM_d0_ivl_869
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2970
  U3127: xor_HPC2
    port map (
      a => LPM_q_ivl_877,
      b => LPM_q_ivl_888,
      c => LPM_d0_ivl_898
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2971
  U3128: xor_HPC2
    port map (
      a => LPM_q_ivl_906,
      b => LPM_q_ivl_917,
      c => LPM_d0_ivl_927
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2972
  U3129: xor_HPC2
    port map (
      a => LPM_q_ivl_935,
      b => LPM_q_ivl_946,
      c => LPM_d0_ivl_956
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2973
  U3130: xor_HPC2
    port map (
      a => LPM_q_ivl_964,
      b => LPM_q_ivl_975,
      c => LPM_d0_ivl_985
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2974
  U3131: xor_HPC2
    port map (
      a => LPM_q_ivl_993,
      b => LPM_q_ivl_1004,
      c => LPM_d0_ivl_1014
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2975
  U3132: xor_HPC2
    port map (
      a => LPM_q_ivl_1022,
      b => LPM_q_ivl_1033,
      c => LPM_d0_ivl_1043
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2976
  U3133: xor_HPC2
    port map (
      a => LPM_q_ivl_1051,
      b => LPM_q_ivl_1062,
      c => LPM_d0_ivl_1072
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2977
  U3134: xor_HPC2
    port map (
      a => LPM_q_ivl_1080,
      b => LPM_q_ivl_1091,
      c => LPM_d0_ivl_1101
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2978
  U3135: xor_HPC2
    port map (
      a => LPM_q_ivl_1109,
      b => LPM_q_ivl_1120,
      c => LPM_d0_ivl_1130
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2979
  U3136: xor_HPC2
    port map (
      a => LPM_q_ivl_1138,
      b => LPM_q_ivl_1149,
      c => LPM_d0_ivl_1159
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2980
  U3137: xor_HPC2
    port map (
      a => LPM_q_ivl_1167,
      b => LPM_q_ivl_1178,
      c => LPM_d0_ivl_1188
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2981
  U3138: xor_HPC2
    port map (
      a => LPM_q_ivl_1196,
      b => LPM_q_ivl_1207,
      c => LPM_d0_ivl_1217
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2982
  U3139: xor_HPC2
    port map (
      a => LPM_q_ivl_1225,
      b => LPM_q_ivl_1236,
      c => LPM_d0_ivl_1246
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2983
  U3140: xor_HPC2
    port map (
      a => LPM_q_ivl_1254,
      b => LPM_q_ivl_1265,
      c => LPM_d0_ivl_1275
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2984
  U3141: xor_HPC2
    port map (
      a => LPM_q_ivl_1283,
      b => LPM_q_ivl_1294,
      c => LPM_d0_ivl_1304
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2985
  U3142: xor_HPC2
    port map (
      a => LPM_q_ivl_1312,
      b => LPM_q_ivl_1323,
      c => LPM_d0_ivl_1333
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2986
  U3143: xor_HPC2
    port map (
      a => LPM_q_ivl_1341,
      b => LPM_q_ivl_1352,
      c => LPM_d0_ivl_1362
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2987
  U3144: xor_HPC2
    port map (
      a => LPM_q_ivl_1370,
      b => LPM_q_ivl_1381,
      c => LPM_d0_ivl_1391
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2988
  U3145: xor_HPC2
    port map (
      a => LPM_q_ivl_1399,
      b => LPM_q_ivl_1410,
      c => LPM_d0_ivl_1420
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2989
  U3146: xor_HPC2
    port map (
      a => LPM_q_ivl_1428,
      b => LPM_q_ivl_1439,
      c => LPM_d0_ivl_1449
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2990
  U3147: xor_HPC2
    port map (
      a => LPM_q_ivl_1457,
      b => LPM_q_ivl_1468,
      c => LPM_d0_ivl_1478
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2991
  U3148: xor_HPC2
    port map (
      a => LPM_q_ivl_1486,
      b => LPM_q_ivl_1497,
      c => LPM_d0_ivl_1507
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2992
  U3149: xor_HPC2
    port map (
      a => LPM_q_ivl_1515,
      b => LPM_q_ivl_1526,
      c => LPM_d0_ivl_1536
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2993
  U3150: xor_HPC2
    port map (
      a => LPM_q_ivl_1544,
      b => LPM_q_ivl_1555,
      c => LPM_d0_ivl_1565
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2994
  U3151: xor_HPC2
    port map (
      a => LPM_q_ivl_1573,
      b => LPM_q_ivl_1584,
      c => LPM_d0_ivl_1594
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2995
  U3152: xor_HPC2
    port map (
      a => LPM_q_ivl_1602,
      b => LPM_q_ivl_1613,
      c => LPM_d0_ivl_1623
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2996
  U3153: xor_HPC2
    port map (
      a => LPM_q_ivl_1631,
      b => LPM_q_ivl_1642,
      c => LPM_d0_ivl_1652
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2997
  U3154: xor_HPC2
    port map (
      a => LPM_q_ivl_1660,
      b => LPM_q_ivl_1671,
      c => LPM_d0_ivl_1681
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2998
  U3155: xor_HPC2
    port map (
      a => LPM_q_ivl_1689,
      b => LPM_q_ivl_1700,
      c => LPM_d0_ivl_1710
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:2999
  U3156: xor_HPC2
    port map (
      a => LPM_q_ivl_1718,
      b => LPM_q_ivl_1729,
      c => LPM_d0_ivl_1739
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3000
  U3157: xor_HPC2
    port map (
      a => LPM_q_ivl_1747,
      b => LPM_q_ivl_1758,
      c => LPM_d0_ivl_1768
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3001
  U3158: xor_HPC2
    port map (
      a => LPM_q_ivl_1776,
      b => LPM_q_ivl_1787,
      c => LPM_d0_ivl_1797
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3002
  U3159: xor_HPC2
    port map (
      a => LPM_q_ivl_1805,
      b => LPM_q_ivl_1816,
      c => LPM_d0_ivl_1826
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3003
  U3160: xor_HPC2
    port map (
      a => LPM_q_ivl_1834,
      b => LPM_q_ivl_1845,
      c => LPM_d0_ivl_1855
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3004
  U3161: xor_HPC2
    port map (
      a => LPM_q_ivl_1863,
      b => LPM_q_ivl_1874,
      c => LPM_d0_ivl_1884
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3005
  U3162: xor_HPC2
    port map (
      a => LPM_q_ivl_1892,
      b => LPM_q_ivl_1903,
      c => LPM_d0_ivl_1913
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3006
  U3163: xor_HPC2
    port map (
      a => LPM_q_ivl_1921,
      b => LPM_q_ivl_1932,
      c => LPM_d0_ivl_1942
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3007
  U3164: xor_HPC2
    port map (
      a => LPM_q_ivl_1950,
      b => LPM_q_ivl_1961,
      c => LPM_d0_ivl_1971
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3008
  U3165: xor_HPC2
    port map (
      a => LPM_q_ivl_1979,
      b => LPM_q_ivl_1990,
      c => LPM_d0_ivl_2000
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3009
  U3166: xor_HPC2
    port map (
      a => LPM_q_ivl_2008,
      b => LPM_q_ivl_2019,
      c => LPM_d0_ivl_2029
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3010
  U3167: xor_HPC2
    port map (
      a => LPM_q_ivl_2037,
      b => LPM_q_ivl_2048,
      c => LPM_d0_ivl_2058
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3011
  U3168: xor_HPC2
    port map (
      a => LPM_q_ivl_2066,
      b => LPM_q_ivl_2077,
      c => LPM_d0_ivl_2087
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3012
  U3169: xor_HPC2
    port map (
      a => LPM_q_ivl_2095,
      b => LPM_q_ivl_2106,
      c => LPM_d0_ivl_2116
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3013
  U3170: xor_HPC2
    port map (
      a => LPM_q_ivl_2124,
      b => LPM_q_ivl_2135,
      c => LPM_d0_ivl_2145
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3014
  U3171: xor_HPC2
    port map (
      a => LPM_q_ivl_2153,
      b => LPM_q_ivl_2164,
      c => LPM_d0_ivl_2174
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3015
  U3172: xor_HPC2
    port map (
      a => LPM_q_ivl_2182,
      b => LPM_q_ivl_2193,
      c => LPM_d0_ivl_2203
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3016
  U3173: xor_HPC2
    port map (
      a => LPM_q_ivl_2211,
      b => LPM_q_ivl_2222,
      c => LPM_d0_ivl_2232
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3017
  U3174: xor_HPC2
    port map (
      a => LPM_q_ivl_2240,
      b => LPM_q_ivl_2251,
      c => LPM_d0_ivl_2261
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3018
  U3175: xor_HPC2
    port map (
      a => LPM_q_ivl_2269,
      b => LPM_q_ivl_2280,
      c => LPM_d0_ivl_2290
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3019
  U3176: xor_HPC2
    port map (
      a => LPM_q_ivl_2298,
      b => LPM_q_ivl_2309,
      c => LPM_d0_ivl_2319
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3020
  U3177: xor_HPC2
    port map (
      a => LPM_q_ivl_2327,
      b => LPM_q_ivl_2338,
      c => LPM_d0_ivl_2348
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3021
  U3178: xor_HPC2
    port map (
      a => LPM_q_ivl_2356,
      b => LPM_q_ivl_2367,
      c => LPM_d0_ivl_2377
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3022
  U3179: xor_HPC2
    port map (
      a => LPM_q_ivl_2385,
      b => LPM_q_ivl_2396,
      c => LPM_d0_ivl_2406
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3023
  U3180: xor_HPC2
    port map (
      a => LPM_q_ivl_2414,
      b => LPM_q_ivl_2425,
      c => LPM_d0_ivl_2435
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3024
  U3181: xor_HPC2
    port map (
      a => LPM_q_ivl_2443,
      b => LPM_q_ivl_2454,
      c => LPM_d0_ivl_2464
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3025
  U3182: xor_HPC2
    port map (
      a => LPM_q_ivl_2472,
      b => LPM_q_ivl_2483,
      c => LPM_d0_ivl_2493
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3026
  U3183: xor_HPC2
    port map (
      a => LPM_q_ivl_2501,
      b => LPM_q_ivl_2512,
      c => LPM_d0_ivl_2522
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3027
  U3184: xor_HPC2
    port map (
      a => LPM_q_ivl_2530,
      b => LPM_q_ivl_2541,
      c => LPM_d0_ivl_2551
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3028
  U3185: xor_HPC2
    port map (
      a => LPM_q_ivl_2559,
      b => LPM_q_ivl_2570,
      c => LPM_d0_ivl_2580
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3029
  U3186: xor_HPC2
    port map (
      a => LPM_q_ivl_2588,
      b => LPM_q_ivl_2599,
      c => LPM_d0_ivl_2609
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3030
  U3187: xor_HPC2
    port map (
      a => LPM_q_ivl_2617,
      b => LPM_q_ivl_2628,
      c => LPM_d0_ivl_2638
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3031
  U3188: xor_HPC2
    port map (
      a => LPM_q_ivl_2646,
      b => LPM_q_ivl_2657,
      c => LPM_d0_ivl_2667
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3032
  U3189: xor_HPC2
    port map (
      a => LPM_q_ivl_2675,
      b => LPM_q_ivl_2686,
      c => LPM_d0_ivl_2696
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3033
  U3190: xor_HPC2
    port map (
      a => LPM_q_ivl_2704,
      b => LPM_q_ivl_2715,
      c => LPM_d0_ivl_2725
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3034
  U3191: xor_HPC2
    port map (
      a => LPM_q_ivl_2733,
      b => LPM_q_ivl_2744,
      c => LPM_d0_ivl_2754
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3035
  U3192: xor_HPC2
    port map (
      a => LPM_q_ivl_2762,
      b => LPM_q_ivl_2773,
      c => LPM_d0_ivl_2783
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3036
  U3193: xor_HPC2
    port map (
      a => LPM_q_ivl_2791,
      b => LPM_q_ivl_2802,
      c => LPM_d0_ivl_2812
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3037
  U3194: xor_HPC2
    port map (
      a => LPM_q_ivl_2820,
      b => LPM_q_ivl_2831,
      c => LPM_d0_ivl_2841
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3038
  U3195: xor_HPC2
    port map (
      a => LPM_q_ivl_2849,
      b => LPM_q_ivl_2860,
      c => LPM_d0_ivl_2870
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3039
  U3196: xor_HPC2
    port map (
      a => LPM_q_ivl_2878,
      b => LPM_q_ivl_2889,
      c => LPM_d0_ivl_2899
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3040
  U3197: xor_HPC2
    port map (
      a => LPM_q_ivl_2907,
      b => LPM_q_ivl_2918,
      c => LPM_d0_ivl_2928
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3041
  U3198: xor_HPC2
    port map (
      a => LPM_q_ivl_2936,
      b => LPM_q_ivl_2947,
      c => LPM_d0_ivl_2957
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3042
  U3199: xor_HPC2
    port map (
      a => LPM_q_ivl_2965,
      b => LPM_q_ivl_2976,
      c => LPM_d0_ivl_2986
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3043
  U3200: xor_HPC2
    port map (
      a => LPM_q_ivl_2994,
      b => LPM_q_ivl_3005,
      c => LPM_d0_ivl_3015
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3044
  U3201: xor_HPC2
    port map (
      a => LPM_q_ivl_3023,
      b => LPM_q_ivl_3034,
      c => LPM_d0_ivl_3044
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3045
  U3202: xor_HPC2
    port map (
      a => LPM_q_ivl_3052,
      b => LPM_q_ivl_3063,
      c => LPM_d0_ivl_3073
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3046
  U3203: xor_HPC2
    port map (
      a => LPM_q_ivl_3081,
      b => LPM_q_ivl_3092,
      c => LPM_d0_ivl_3102
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3047
  U3204: xor_HPC2
    port map (
      a => LPM_q_ivl_3110,
      b => LPM_q_ivl_3121,
      c => LPM_d0_ivl_3131
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3048
  U3205: xor_HPC2
    port map (
      a => LPM_q_ivl_3139,
      b => LPM_q_ivl_3150,
      c => LPM_d0_ivl_3160
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3049
  U3206: xor_HPC2
    port map (
      a => LPM_q_ivl_3168,
      b => LPM_q_ivl_3179,
      c => LPM_d0_ivl_3189
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3050
  U3207: xor_HPC2
    port map (
      a => LPM_q_ivl_3197,
      b => LPM_q_ivl_3208,
      c => LPM_d0_ivl_3218
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3051
  U3208: xor_HPC2
    port map (
      a => LPM_q_ivl_3226,
      b => LPM_q_ivl_3237,
      c => LPM_d0_ivl_3247
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3052
  U3209: xor_HPC2
    port map (
      a => LPM_q_ivl_3255,
      b => LPM_q_ivl_3266,
      c => LPM_d0_ivl_3276
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3053
  U3210: xor_HPC2
    port map (
      a => LPM_q_ivl_3284,
      b => LPM_q_ivl_3295,
      c => LPM_d0_ivl_3305
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3054
  U3211: xor_HPC2
    port map (
      a => LPM_q_ivl_3313,
      b => LPM_q_ivl_3324,
      c => LPM_d0_ivl_3334
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3055
  U3212: xor_HPC2
    port map (
      a => LPM_q_ivl_3342,
      b => LPM_q_ivl_3353,
      c => LPM_d0_ivl_3363
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3056
  U3213: xor_HPC2
    port map (
      a => LPM_q_ivl_3371,
      b => LPM_q_ivl_3382,
      c => LPM_d0_ivl_3392
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3057
  U3214: xor_HPC2
    port map (
      a => LPM_q_ivl_3400,
      b => LPM_q_ivl_3411,
      c => LPM_d0_ivl_3421
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3058
  U3215: xor_HPC2
    port map (
      a => LPM_q_ivl_3429,
      b => LPM_q_ivl_3440,
      c => LPM_d0_ivl_3450
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3059
  U3216: xor_HPC2
    port map (
      a => LPM_q_ivl_3458,
      b => LPM_q_ivl_3469,
      c => LPM_d0_ivl_3479
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3060
  U3217: xor_HPC2
    port map (
      a => LPM_q_ivl_3487,
      b => LPM_q_ivl_3498,
      c => LPM_d0_ivl_3508
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3061
  U3218: xor_HPC2
    port map (
      a => LPM_q_ivl_3516,
      b => LPM_q_ivl_3527,
      c => LPM_d0_ivl_3537
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3062
  U3219: xor_HPC2
    port map (
      a => LPM_q_ivl_3545,
      b => LPM_q_ivl_3556,
      c => LPM_d0_ivl_3566
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3063
  U3220: xor_HPC2
    port map (
      a => LPM_q_ivl_3574,
      b => LPM_q_ivl_3585,
      c => LPM_d0_ivl_3595
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3064
  U3221: xor_HPC2
    port map (
      a => LPM_q_ivl_3603,
      b => LPM_q_ivl_3614,
      c => LPM_d0_ivl_3624
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3065
  U3222: xor_HPC2
    port map (
      a => LPM_q_ivl_3632,
      b => LPM_q_ivl_3643,
      c => LPM_d0_ivl_3653
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3066
  U3223: xor_HPC2
    port map (
      a => LPM_q_ivl_3661,
      b => LPM_q_ivl_3672,
      c => LPM_d0_ivl_3682
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3067
  U3224: xor_HPC2
    port map (
      a => LPM_q_ivl_3690,
      b => LPM_q_ivl_3701,
      c => LPM_d0_ivl_3711
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3361
  U3225: xnor_HPC2
    port map (
      a => LPM_q_ivl_7692,
      b => LPM_q_ivl_7701,
      c => LPM_d0_ivl_7709
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3362
  U3226: xnor_HPC2
    port map (
      a => LPM_q_ivl_7717,
      b => LPM_q_ivl_7724,
      c => LPM_d0_ivl_7732
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3363
  U3227: xnor_HPC2
    port map (
      a => LPM_q_ivl_7740,
      b => LPM_q_ivl_7749,
      c => LPM_d0_ivl_7757
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3364
  U3228: xnor_HPC2
    port map (
      a => LPM_q_ivl_7765,
      b => LPM_q_ivl_7772,
      c => LPM_d0_ivl_7780
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3365
  U3229: xnor_HPC2
    port map (
      a => LPM_q_ivl_7784,
      b => LPM_q_ivl_7791,
      c => LPM_d0_ivl_7799
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3366
  U3230: xnor_HPC2
    port map (
      a => LPM_q_ivl_7807,
      b => LPM_q_ivl_7816,
      c => LPM_d0_ivl_7824
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3367
  U3231: xnor_HPC2
    port map (
      a => LPM_q_ivl_7832,
      b => LPM_q_ivl_7839,
      c => LPM_d0_ivl_7847
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3368
  U3232: xnor_HPC2
    port map (
      a => LPM_q_ivl_7851,
      b => LPM_q_ivl_7858,
      c => LPM_d0_ivl_7870
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3369
  U3233: xnor_HPC2
    port map (
      a => LPM_q_ivl_7878,
      b => LPM_q_ivl_7887,
      c => LPM_d0_ivl_7895
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3370
  U3234: xnor_HPC2
    port map (
      a => LPM_q_ivl_7903,
      b => LPM_q_ivl_7910,
      c => LPM_d0_ivl_7918
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3371
  U3235: xnor_HPC2
    port map (
      a => LPM_q_ivl_7926,
      b => LPM_q_ivl_7935,
      c => LPM_d0_ivl_7943
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3372
  U3236: xnor_HPC2
    port map (
      a => LPM_q_ivl_7951,
      b => LPM_q_ivl_7958,
      c => LPM_d0_ivl_7966
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3373
  U3237: xnor_HPC2
    port map (
      a => LPM_q_ivl_7970,
      b => LPM_q_ivl_7977,
      c => LPM_d0_ivl_7985
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3374
  U3238: xnor_HPC2
    port map (
      a => LPM_q_ivl_7993,
      b => LPM_q_ivl_8002,
      c => LPM_d0_ivl_8010
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3375
  U3239: xnor_HPC2
    port map (
      a => LPM_q_ivl_8018,
      b => LPM_q_ivl_8025,
      c => LPM_d0_ivl_8033
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3376
  U3240: xnor_HPC2
    port map (
      a => LPM_q_ivl_8037,
      b => LPM_q_ivl_8044,
      c => LPM_d0_ivl_8056
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3377
  U3241: xnor_HPC2
    port map (
      a => LPM_q_ivl_8064,
      b => LPM_q_ivl_8073,
      c => LPM_d0_ivl_8081
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3378
  U3242: xnor_HPC2
    port map (
      a => LPM_q_ivl_8089,
      b => LPM_q_ivl_8096,
      c => LPM_d0_ivl_8104
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3379
  U3243: xnor_HPC2
    port map (
      a => LPM_q_ivl_8112,
      b => LPM_q_ivl_8121,
      c => LPM_d0_ivl_8129
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3380
  U3244: xnor_HPC2
    port map (
      a => LPM_q_ivl_8137,
      b => LPM_q_ivl_8144,
      c => LPM_d0_ivl_8152
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3381
  U3245: xnor_HPC2
    port map (
      a => LPM_q_ivl_8156,
      b => LPM_q_ivl_8163,
      c => LPM_d0_ivl_8171
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3382
  U3246: xnor_HPC2
    port map (
      a => LPM_q_ivl_8179,
      b => LPM_q_ivl_8188,
      c => LPM_d0_ivl_8196
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3383
  U3247: xnor_HPC2
    port map (
      a => LPM_q_ivl_8204,
      b => LPM_q_ivl_8211,
      c => LPM_d0_ivl_8219
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3384
  U3248: xnor_HPC2
    port map (
      a => LPM_q_ivl_8223,
      b => LPM_q_ivl_8230,
      c => LPM_d0_ivl_8242
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3385
  U3249: xnor_HPC2
    port map (
      a => LPM_q_ivl_8250,
      b => LPM_q_ivl_8259,
      c => LPM_d0_ivl_8267
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3386
  U3250: xnor_HPC2
    port map (
      a => LPM_q_ivl_8275,
      b => LPM_q_ivl_8282,
      c => LPM_d0_ivl_8290
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3387
  U3251: xnor_HPC2
    port map (
      a => LPM_q_ivl_8298,
      b => LPM_q_ivl_8307,
      c => LPM_d0_ivl_8315
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3388
  U3252: xnor_HPC2
    port map (
      a => LPM_q_ivl_8323,
      b => LPM_q_ivl_8330,
      c => LPM_d0_ivl_8338
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3389
  U3253: xnor_HPC2
    port map (
      a => LPM_q_ivl_8342,
      b => LPM_q_ivl_8349,
      c => LPM_d0_ivl_8357
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3390
  U3254: xnor_HPC2
    port map (
      a => LPM_q_ivl_8365,
      b => LPM_q_ivl_8374,
      c => LPM_d0_ivl_8382
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3391
  U3255: xnor_HPC2
    port map (
      a => LPM_q_ivl_8390,
      b => LPM_q_ivl_8397,
      c => LPM_d0_ivl_8405
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3392
  U3256: xnor_HPC2
    port map (
      a => LPM_q_ivl_8409,
      b => LPM_q_ivl_8416,
      c => LPM_d0_ivl_8428
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3393
  U3257: xnor_HPC2
    port map (
      a => LPM_q_ivl_8436,
      b => LPM_q_ivl_8445,
      c => LPM_d0_ivl_8453
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3394
  U3258: xnor_HPC2
    port map (
      a => LPM_q_ivl_8461,
      b => LPM_q_ivl_8468,
      c => LPM_d0_ivl_8476
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3395
  U3259: xnor_HPC2
    port map (
      a => LPM_q_ivl_8484,
      b => LPM_q_ivl_8493,
      c => LPM_d0_ivl_8501
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3396
  U3260: xnor_HPC2
    port map (
      a => LPM_q_ivl_8509,
      b => LPM_q_ivl_8516,
      c => LPM_d0_ivl_8524
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3397
  U3261: xnor_HPC2
    port map (
      a => LPM_q_ivl_8528,
      b => LPM_q_ivl_8535,
      c => LPM_d0_ivl_8543
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3398
  U3262: xnor_HPC2
    port map (
      a => LPM_q_ivl_8551,
      b => LPM_q_ivl_8560,
      c => LPM_d0_ivl_8568
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3399
  U3263: xnor_HPC2
    port map (
      a => LPM_q_ivl_8576,
      b => LPM_q_ivl_8583,
      c => LPM_d0_ivl_8591
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3400
  U3264: xnor_HPC2
    port map (
      a => LPM_q_ivl_8595,
      b => LPM_q_ivl_8602,
      c => LPM_d0_ivl_8614
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3401
  U3265: xnor_HPC2
    port map (
      a => LPM_q_ivl_8622,
      b => LPM_q_ivl_8631,
      c => LPM_d0_ivl_8639
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3402
  U3266: xnor_HPC2
    port map (
      a => LPM_q_ivl_8647,
      b => LPM_q_ivl_8654,
      c => LPM_d0_ivl_8662
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3403
  U3267: xnor_HPC2
    port map (
      a => LPM_q_ivl_8670,
      b => LPM_q_ivl_8679,
      c => LPM_d0_ivl_8687
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3404
  U3268: xnor_HPC2
    port map (
      a => LPM_q_ivl_8695,
      b => LPM_q_ivl_8702,
      c => LPM_d0_ivl_8710
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3405
  U3269: xnor_HPC2
    port map (
      a => LPM_q_ivl_8714,
      b => LPM_q_ivl_8721,
      c => LPM_d0_ivl_8729
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3406
  U3270: xnor_HPC2
    port map (
      a => LPM_q_ivl_8737,
      b => LPM_q_ivl_8746,
      c => LPM_d0_ivl_8754
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3407
  U3271: xnor_HPC2
    port map (
      a => LPM_q_ivl_8762,
      b => LPM_q_ivl_8769,
      c => LPM_d0_ivl_8777
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3408
  U3272: xnor_HPC2
    port map (
      a => LPM_q_ivl_8781,
      b => LPM_q_ivl_8788,
      c => LPM_d0_ivl_8800
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3409
  U3273: xnor_HPC2
    port map (
      a => LPM_q_ivl_8808,
      b => LPM_q_ivl_8817,
      c => LPM_d0_ivl_8825
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3410
  U3274: xnor_HPC2
    port map (
      a => LPM_q_ivl_8833,
      b => LPM_q_ivl_8840,
      c => LPM_d0_ivl_8848
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3411
  U3275: xnor_HPC2
    port map (
      a => LPM_q_ivl_8852,
      b => LPM_q_ivl_8859,
      c => LPM_d0_ivl_8867
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3412
  U3276: xnor_HPC2
    port map (
      a => LPM_q_ivl_8875,
      b => LPM_q_ivl_8884,
      c => LPM_d0_ivl_8892
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3413
  U3277: xnor_HPC2
    port map (
      a => LPM_q_ivl_8900,
      b => LPM_q_ivl_8907,
      c => LPM_d0_ivl_8915
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3414
  U3278: xnor_HPC2
    port map (
      a => LPM_q_ivl_8919,
      b => LPM_q_ivl_8926,
      c => LPM_d0_ivl_8938
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3415
  U3279: xnor_HPC2
    port map (
      a => LPM_q_ivl_8946,
      b => LPM_q_ivl_8955,
      c => LPM_d0_ivl_8963
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3416
  U3280: xnor_HPC2
    port map (
      a => LPM_q_ivl_8971,
      b => LPM_q_ivl_8978,
      c => LPM_d0_ivl_8986
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3417
  U3281: xnor_HPC2
    port map (
      a => LPM_q_ivl_8994,
      b => LPM_q_ivl_9003,
      c => LPM_d0_ivl_9011
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3418
  U3282: xnor_HPC2
    port map (
      a => LPM_q_ivl_9019,
      b => LPM_q_ivl_9026,
      c => LPM_d0_ivl_9034
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3419
  U3283: xnor_HPC2
    port map (
      a => LPM_q_ivl_9038,
      b => LPM_q_ivl_9045,
      c => LPM_d0_ivl_9053
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3420
  U3284: xnor_HPC2
    port map (
      a => LPM_q_ivl_9061,
      b => LPM_q_ivl_9070,
      c => LPM_d0_ivl_9078
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3421
  U3285: xnor_HPC2
    port map (
      a => LPM_q_ivl_9086,
      b => LPM_q_ivl_9093,
      c => LPM_d0_ivl_9101
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3422
  U3286: xnor_HPC2
    port map (
      a => LPM_q_ivl_9105,
      b => LPM_q_ivl_9112,
      c => LPM_d0_ivl_9124
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3423
  U3287: xnor_HPC2
    port map (
      a => LPM_q_ivl_9132,
      b => LPM_q_ivl_9141,
      c => LPM_d0_ivl_9149
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3424
  U3288: xnor_HPC2
    port map (
      a => LPM_q_ivl_9157,
      b => LPM_q_ivl_9164,
      c => LPM_d0_ivl_9172
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3425
  U3289: xnor_HPC2
    port map (
      a => LPM_q_ivl_9176,
      b => LPM_q_ivl_9183,
      c => LPM_d0_ivl_9191
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3426
  U3290: xnor_HPC2
    port map (
      a => LPM_q_ivl_9199,
      b => LPM_q_ivl_9208,
      c => LPM_d0_ivl_9216
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3427
  U3291: xnor_HPC2
    port map (
      a => LPM_q_ivl_9224,
      b => LPM_q_ivl_9231,
      c => LPM_d0_ivl_9239
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3428
  U3292: xnor_HPC2
    port map (
      a => LPM_q_ivl_9243,
      b => LPM_q_ivl_9250,
      c => LPM_d0_ivl_9262
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3429
  U3293: xnor_HPC2
    port map (
      a => LPM_q_ivl_9270,
      b => LPM_q_ivl_9279,
      c => LPM_d0_ivl_9287
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3430
  U3294: xnor_HPC2
    port map (
      a => LPM_q_ivl_9295,
      b => LPM_q_ivl_9302,
      c => LPM_d0_ivl_9310
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3431
  U3295: xnor_HPC2
    port map (
      a => LPM_q_ivl_9314,
      b => LPM_q_ivl_9321,
      c => LPM_d0_ivl_9329
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3432
  U3296: xnor_HPC2
    port map (
      a => LPM_q_ivl_9337,
      b => LPM_q_ivl_9346,
      c => LPM_d0_ivl_9354
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3433
  U3297: xnor_HPC2
    port map (
      a => LPM_q_ivl_9362,
      b => LPM_q_ivl_9369,
      c => LPM_d0_ivl_9377
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3434
  U3298: xnor_HPC2
    port map (
      a => LPM_q_ivl_9381,
      b => LPM_q_ivl_9388,
      c => LPM_d0_ivl_9400
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3435
  U3299: xnor_HPC2
    port map (
      a => LPM_q_ivl_9408,
      b => LPM_q_ivl_9417,
      c => LPM_d0_ivl_9425
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3436
  U3300: xnor_HPC2
    port map (
      a => LPM_q_ivl_9433,
      b => LPM_q_ivl_9440,
      c => LPM_d0_ivl_9448
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3437
  U3301: xnor_HPC2
    port map (
      a => LPM_q_ivl_9452,
      b => LPM_q_ivl_9459,
      c => LPM_d0_ivl_9467
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3438
  U3302: xnor_HPC2
    port map (
      a => LPM_q_ivl_9475,
      b => LPM_q_ivl_9484,
      c => LPM_d0_ivl_9492
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3439
  U3303: xnor_HPC2
    port map (
      a => LPM_q_ivl_9500,
      b => LPM_q_ivl_9507,
      c => LPM_d0_ivl_9515
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3440
  U3304: xnor_HPC2
    port map (
      a => LPM_q_ivl_9519,
      b => LPM_q_ivl_9526,
      c => LPM_d0_ivl_9538
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3441
  U3305: xnor_HPC2
    port map (
      a => LPM_q_ivl_9546,
      b => LPM_q_ivl_9555,
      c => LPM_d0_ivl_9563
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3442
  U3306: xnor_HPC2
    port map (
      a => LPM_q_ivl_9571,
      b => LPM_q_ivl_9578,
      c => LPM_d0_ivl_9586
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3443
  U3307: xnor_HPC2
    port map (
      a => LPM_q_ivl_9590,
      b => LPM_q_ivl_9597,
      c => LPM_d0_ivl_9605
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3444
  U3308: xnor_HPC2
    port map (
      a => LPM_q_ivl_9613,
      b => LPM_q_ivl_9622,
      c => LPM_d0_ivl_9630
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3445
  U3309: xnor_HPC2
    port map (
      a => LPM_q_ivl_9638,
      b => LPM_q_ivl_9645,
      c => LPM_d0_ivl_9653
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3446
  U3310: xnor_HPC2
    port map (
      a => LPM_q_ivl_9657,
      b => LPM_q_ivl_9664,
      c => LPM_d0_ivl_9676
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3447
  U3311: xnor_HPC2
    port map (
      a => LPM_q_ivl_9680,
      b => LPM_q_ivl_9687,
      c => LPM_d0_ivl_9695
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3448
  U3312: xnor_HPC2
    port map (
      a => LPM_q_ivl_9703,
      b => LPM_q_ivl_9712,
      c => LPM_d0_ivl_9720
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3449
  U3313: xnor_HPC2
    port map (
      a => LPM_q_ivl_9728,
      b => LPM_q_ivl_9735,
      c => LPM_d0_ivl_9743
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3450
  U3314: xnor_HPC2
    port map (
      a => LPM_q_ivl_9747,
      b => LPM_q_ivl_9754,
      c => LPM_d0_ivl_9766
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3451
  U3315: xnor_HPC2
    port map (
      a => LPM_q_ivl_9770,
      b => LPM_q_ivl_9777,
      c => LPM_d0_ivl_9785
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3452
  U3316: xnor_HPC2
    port map (
      a => LPM_q_ivl_9793,
      b => LPM_q_ivl_9802,
      c => LPM_d0_ivl_9810
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3453
  U3317: xnor_HPC2
    port map (
      a => LPM_q_ivl_9818,
      b => LPM_q_ivl_9825,
      c => LPM_d0_ivl_9833
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3454
  U3318: xnor_HPC2
    port map (
      a => LPM_q_ivl_9837,
      b => LPM_q_ivl_9844,
      c => LPM_d0_ivl_9856
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3455
  U3319: xnor_HPC2
    port map (
      a => LPM_q_ivl_9864,
      b => LPM_q_ivl_9873,
      c => LPM_d0_ivl_9881
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3456
  U3320: xnor_HPC2
    port map (
      a => LPM_q_ivl_9889,
      b => LPM_q_ivl_9896,
      c => LPM_d0_ivl_9904
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3457
  U3321: xnor_HPC2
    port map (
      a => LPM_q_ivl_9908,
      b => LPM_q_ivl_9915,
      c => LPM_d0_ivl_9923
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3458
  U3322: xnor_HPC2
    port map (
      a => LPM_q_ivl_9931,
      b => LPM_q_ivl_9940,
      c => LPM_d0_ivl_9948
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3459
  U3323: xnor_HPC2
    port map (
      a => LPM_q_ivl_9956,
      b => LPM_q_ivl_9963,
      c => LPM_d0_ivl_9971
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3460
  U3324: xnor_HPC2
    port map (
      a => LPM_q_ivl_9975,
      b => LPM_q_ivl_9982,
      c => LPM_d0_ivl_9994
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3461
  U3325: xnor_HPC2
    port map (
      a => LPM_q_ivl_10002,
      b => LPM_q_ivl_10011,
      c => LPM_d0_ivl_10019
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3462
  U3326: xnor_HPC2
    port map (
      a => LPM_q_ivl_10027,
      b => LPM_q_ivl_10034,
      c => LPM_d0_ivl_10042
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3463
  U3327: xnor_HPC2
    port map (
      a => LPM_q_ivl_10046,
      b => LPM_q_ivl_10053,
      c => LPM_d0_ivl_10061
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3464
  U3328: xnor_HPC2
    port map (
      a => LPM_q_ivl_10069,
      b => LPM_q_ivl_10078,
      c => LPM_d0_ivl_10086
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3465
  U3329: xnor_HPC2
    port map (
      a => LPM_q_ivl_10094,
      b => LPM_q_ivl_10101,
      c => LPM_d0_ivl_10109
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3466
  U3330: xnor_HPC2
    port map (
      a => LPM_q_ivl_10113,
      b => LPM_q_ivl_10120,
      c => LPM_d0_ivl_10132
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3467
  U3331: xor_HPC2
    port map (
      a => LPM_q_ivl_10138,
      b => LPM_q_ivl_10149,
      c => LPM_d0_ivl_10157
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3468
  U3332: xor_HPC2
    port map (
      a => LPM_q_ivl_10163,
      b => LPM_q_ivl_10170,
      c => LPM_d0_ivl_10178
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3068
  U3333: xnor_HPC2
    port map (
      a => LPM_q_ivl_3719,
      b => LPM_q_ivl_3730,
      c => LPM_d0_ivl_3738
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3469
  U3334: xnor_HPC2
    port map (
      a => LPM_q_ivl_10182,
      b => LPM_q_ivl_10189,
      c => LPM_d0_ivl_10197
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3470
  U3335: xor_HPC2
    port map (
      a => LPM_q_ivl_10203,
      b => LPM_q_ivl_10214,
      c => LPM_d0_ivl_10222
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3471
  U3336: xor_HPC2
    port map (
      a => LPM_q_ivl_10228,
      b => LPM_q_ivl_10239,
      c => LPM_d0_ivl_10247
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3472
  U3337: xnor_HPC2
    port map (
      a => LPM_q_ivl_10255,
      b => LPM_q_ivl_10262,
      c => LPM_d0_ivl_10270
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3473
  U3338: xnor_HPC2
    port map (
      a => LPM_q_ivl_10274,
      b => LPM_q_ivl_10281,
      c => LPM_d0_ivl_10289
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3474
  U3339: xnor_HPC2
    port map (
      a => LPM_q_ivl_10293,
      b => LPM_q_ivl_10300,
      c => LPM_d0_ivl_10308
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3475
  U3340: xor_HPC2
    port map (
      a => LPM_q_ivl_10314,
      b => LPM_q_ivl_10325,
      c => LPM_d0_ivl_10333
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3476
  U3341: xor_HPC2
    port map (
      a => LPM_q_ivl_10339,
      b => LPM_q_ivl_10350,
      c => LPM_d0_ivl_10358
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3477
  U3342: xnor_HPC2
    port map (
      a => LPM_q_ivl_10366,
      b => LPM_q_ivl_10373,
      c => LPM_d0_ivl_10381
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3478
  U3343: xnor_HPC2
    port map (
      a => LPM_q_ivl_10385,
      b => LPM_q_ivl_10392,
      c => LPM_d0_ivl_10400
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3479
  U3344: xnor_HPC2
    port map (
      a => LPM_q_ivl_10404,
      b => LPM_q_ivl_10411,
      c => LPM_d0_ivl_10423
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3480
  U3345: xor_HPC2
    port map (
      a => LPM_q_ivl_10429,
      b => LPM_q_ivl_10440,
      c => LPM_d0_ivl_10448
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3481
  U3346: xor_HPC2
    port map (
      a => LPM_q_ivl_10454,
      b => LPM_q_ivl_10461,
      c => LPM_d0_ivl_10469
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3069
  U3347: xnor_HPC2
    port map (
      a => LPM_q_ivl_3746,
      b => LPM_q_ivl_3757,
      c => LPM_d0_ivl_3765
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3482
  U3348: xnor_HPC2
    port map (
      a => LPM_q_ivl_10473,
      b => LPM_q_ivl_10480,
      c => LPM_d0_ivl_10488
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3483
  U3349: xor_HPC2
    port map (
      a => LPM_q_ivl_10494,
      b => LPM_q_ivl_10505,
      c => LPM_d0_ivl_10513
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3484
  U3350: xor_HPC2
    port map (
      a => LPM_q_ivl_10519,
      b => LPM_q_ivl_10530,
      c => LPM_d0_ivl_10538
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3485
  U3351: xnor_HPC2
    port map (
      a => LPM_q_ivl_10546,
      b => LPM_q_ivl_10553,
      c => LPM_d0_ivl_10561
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3486
  U3352: xnor_HPC2
    port map (
      a => LPM_q_ivl_10565,
      b => LPM_q_ivl_10572,
      c => LPM_d0_ivl_10580
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3487
  U3353: xnor_HPC2
    port map (
      a => LPM_q_ivl_10584,
      b => LPM_q_ivl_10591,
      c => LPM_d0_ivl_10599
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3488
  U3354: xor_HPC2
    port map (
      a => LPM_q_ivl_10605,
      b => LPM_q_ivl_10616,
      c => LPM_d0_ivl_10624
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3489
  U3355: xor_HPC2
    port map (
      a => LPM_q_ivl_10630,
      b => LPM_q_ivl_10641,
      c => LPM_d0_ivl_10649
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3490
  U3356: xnor_HPC2
    port map (
      a => LPM_q_ivl_10657,
      b => LPM_q_ivl_10664,
      c => LPM_d0_ivl_10672
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3491
  U3357: xnor_HPC2
    port map (
      a => LPM_q_ivl_10676,
      b => LPM_q_ivl_10683,
      c => LPM_d0_ivl_10691
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3492
  U3358: xnor_HPC2
    port map (
      a => LPM_q_ivl_10695,
      b => LPM_q_ivl_10702,
      c => LPM_d0_ivl_10714
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3493
  U3359: xnor_HPC2
    port map (
      a => LPM_q_ivl_10718,
      b => LPM_q_ivl_10725,
      c => LPM_d0_ivl_10733
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3494
  U3360: xnor_HPC2
    port map (
      a => LPM_q_ivl_10741,
      b => LPM_q_ivl_10750,
      c => LPM_d0_ivl_10758
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3495
  U3361: xnor_HPC2
    port map (
      a => LPM_q_ivl_10766,
      b => LPM_q_ivl_10773,
      c => LPM_d0_ivl_10781
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3496
  U3362: xnor_HPC2
    port map (
      a => LPM_q_ivl_10785,
      b => LPM_q_ivl_10792,
      c => LPM_d0_ivl_10804
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3497
  U3363: xnor_HPC2
    port map (
      a => LPM_q_ivl_10808,
      b => LPM_q_ivl_10815,
      c => LPM_d0_ivl_10823
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3498
  U3364: xnor_HPC2
    port map (
      a => LPM_q_ivl_10831,
      b => LPM_q_ivl_10840,
      c => LPM_d0_ivl_10848
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3499
  U3365: xnor_HPC2
    port map (
      a => LPM_q_ivl_10856,
      b => LPM_q_ivl_10863,
      c => LPM_d0_ivl_10871
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3500
  U3366: xnor_HPC2
    port map (
      a => LPM_q_ivl_10875,
      b => LPM_q_ivl_10882,
      c => LPM_d0_ivl_10894
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3501
  U3367: xnor_HPC2
    port map (
      a => LPM_q_ivl_10902,
      b => LPM_q_ivl_10911,
      c => LPM_d0_ivl_10919
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3502
  U3368: xnor_HPC2
    port map (
      a => LPM_q_ivl_10927,
      b => LPM_q_ivl_10934,
      c => LPM_d0_ivl_10942
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3503
  U3369: xnor_HPC2
    port map (
      a => LPM_q_ivl_10946,
      b => LPM_q_ivl_10953,
      c => LPM_d0_ivl_10961
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3504
  U3370: xnor_HPC2
    port map (
      a => LPM_q_ivl_10969,
      b => LPM_q_ivl_10978,
      c => LPM_d0_ivl_10986
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3505
  U3371: xnor_HPC2
    port map (
      a => LPM_q_ivl_10994,
      b => LPM_q_ivl_11001,
      c => LPM_d0_ivl_11009
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3506
  U3372: xnor_HPC2
    port map (
      a => LPM_q_ivl_11013,
      b => LPM_q_ivl_11020,
      c => LPM_d0_ivl_11032
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3507
  U3373: xor_HPC2
    port map (
      a => LPM_q_ivl_11038,
      b => LPM_q_ivl_11049,
      c => LPM_d0_ivl_11057
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3508
  U3374: xor_HPC2
    port map (
      a => LPM_q_ivl_11063,
      b => LPM_q_ivl_11074,
      c => LPM_d0_ivl_11082
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3509
  U3375: xnor_HPC2
    port map (
      a => LPM_q_ivl_11090,
      b => LPM_q_ivl_11097,
      c => LPM_d0_ivl_11105
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3510
  U3376: xnor_HPC2
    port map (
      a => LPM_q_ivl_11109,
      b => LPM_q_ivl_11116,
      c => LPM_d0_ivl_11124
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3511
  U3377: xor_HPC2
    port map (
      a => LPM_q_ivl_11130,
      b => LPM_q_ivl_11141,
      c => LPM_d0_ivl_11149
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3512
  U3378: xor_HPC2
    port map (
      a => LPM_q_ivl_11155,
      b => LPM_q_ivl_11162,
      c => LPM_d0_ivl_11170
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3070
  U3379: xnor_HPC2
    port map (
      a => LPM_q_ivl_3773,
      b => LPM_q_ivl_3784,
      c => LPM_d0_ivl_3792
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3513
  U3380: xnor_HPC2
    port map (
      a => LPM_q_ivl_11174,
      b => LPM_q_ivl_11181,
      c => LPM_d0_ivl_11189
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3514
  U3381: xnor_HPC2
    port map (
      a => LPM_q_ivl_11193,
      b => LPM_q_ivl_11200,
      c => LPM_d0_ivl_11208
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3515
  U3382: xor_HPC2
    port map (
      a => LPM_q_ivl_11214,
      b => LPM_q_ivl_11225,
      c => LPM_d0_ivl_11233
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3516
  U3383: xor_HPC2
    port map (
      a => LPM_q_ivl_11239,
      b => LPM_q_ivl_11250,
      c => LPM_d0_ivl_11258
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3517
  U3384: xnor_HPC2
    port map (
      a => LPM_q_ivl_11266,
      b => LPM_q_ivl_11273,
      c => LPM_d0_ivl_11281
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3518
  U3385: xnor_HPC2
    port map (
      a => LPM_q_ivl_11285,
      b => LPM_q_ivl_11292,
      c => LPM_d0_ivl_11300
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3519
  U3386: xnor_HPC2
    port map (
      a => LPM_q_ivl_11304,
      b => LPM_q_ivl_11311,
      c => LPM_d0_ivl_11323
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3520
  U3387: xor_HPC2
    port map (
      a => LPM_q_ivl_11329,
      b => LPM_q_ivl_11340,
      c => LPM_d0_ivl_11348
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3521
  U3388: xor_HPC2
    port map (
      a => LPM_q_ivl_11354,
      b => LPM_q_ivl_11365,
      c => LPM_d0_ivl_11373
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3522
  U3389: xnor_HPC2
    port map (
      a => LPM_q_ivl_11381,
      b => LPM_q_ivl_11388,
      c => LPM_d0_ivl_11396
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3523
  U3390: xnor_HPC2
    port map (
      a => LPM_q_ivl_11400,
      b => LPM_q_ivl_11407,
      c => LPM_d0_ivl_11415
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3524
  U3391: xnor_HPC2
    port map (
      a => LPM_q_ivl_11419,
      b => LPM_q_ivl_11426,
      c => LPM_d0_ivl_11434
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3525
  U3392: xor_HPC2
    port map (
      a => LPM_q_ivl_11440,
      b => LPM_q_ivl_11451,
      c => LPM_d0_ivl_11459
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3526
  U3393: xor_HPC2
    port map (
      a => LPM_q_ivl_11465,
      b => LPM_q_ivl_11472,
      c => LPM_d0_ivl_11480
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3071
  U3394: xnor_HPC2
    port map (
      a => LPM_q_ivl_3800,
      b => LPM_q_ivl_3811,
      c => LPM_d0_ivl_3819
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3527
  U3395: xnor_HPC2
    port map (
      a => LPM_q_ivl_11484,
      b => LPM_q_ivl_11491,
      c => LPM_d0_ivl_11499
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3528
  U3396: xnor_HPC2
    port map (
      a => LPM_q_ivl_11503,
      b => LPM_q_ivl_11510,
      c => LPM_d0_ivl_11522
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3529
  U3397: xor_HPC2
    port map (
      a => LPM_q_ivl_11528,
      b => LPM_q_ivl_11539,
      c => LPM_d0_ivl_11547
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3530
  U3398: xor_HPC2
    port map (
      a => LPM_q_ivl_11553,
      b => LPM_q_ivl_11564,
      c => LPM_d0_ivl_11572
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3531
  U3399: xnor_HPC2
    port map (
      a => LPM_q_ivl_11580,
      b => LPM_q_ivl_11587,
      c => LPM_d0_ivl_11595
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3532
  U3400: xnor_HPC2
    port map (
      a => LPM_q_ivl_11599,
      b => LPM_q_ivl_11606,
      c => LPM_d0_ivl_11614
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3533
  U3401: xnor_HPC2
    port map (
      a => LPM_q_ivl_11618,
      b => LPM_q_ivl_11625,
      c => LPM_d0_ivl_11633
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3534
  U3402: xor_HPC2
    port map (
      a => LPM_q_ivl_11639,
      b => LPM_q_ivl_11650,
      c => LPM_d0_ivl_11658
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3535
  U3403: xor_HPC2
    port map (
      a => LPM_q_ivl_11664,
      b => LPM_q_ivl_11675,
      c => LPM_d0_ivl_11683
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3536
  U3404: xnor_HPC2
    port map (
      a => LPM_q_ivl_11691,
      b => LPM_q_ivl_11698,
      c => LPM_d0_ivl_11706
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3537
  U3405: xnor_HPC2
    port map (
      a => LPM_q_ivl_11710,
      b => LPM_q_ivl_11717,
      c => LPM_d0_ivl_11725
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3538
  U3406: xnor_HPC2
    port map (
      a => LPM_q_ivl_11729,
      b => LPM_q_ivl_11736,
      c => LPM_d0_ivl_11748
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3539
  U3407: xnor_HPC2
    port map (
      a => LPM_q_ivl_11752,
      b => LPM_q_ivl_11759,
      c => LPM_d0_ivl_11767
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3540
  U3408: xnor_HPC2
    port map (
      a => LPM_q_ivl_11775,
      b => LPM_q_ivl_11784,
      c => LPM_d0_ivl_11792
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3541
  U3409: xnor_HPC2
    port map (
      a => LPM_q_ivl_11800,
      b => LPM_q_ivl_11807,
      c => LPM_d0_ivl_11815
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3542
  U3410: xnor_HPC2
    port map (
      a => LPM_q_ivl_11819,
      b => LPM_q_ivl_11826,
      c => LPM_d0_ivl_11838
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3543
  U3411: xnor_HPC2
    port map (
      a => LPM_q_ivl_11842,
      b => LPM_q_ivl_11849,
      c => LPM_d0_ivl_11857
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3544
  U3412: xnor_HPC2
    port map (
      a => LPM_q_ivl_11861,
      b => LPM_q_ivl_11868,
      c => LPM_d0_ivl_11880
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3545
  U3413: xor_HPC2
    port map (
      a => LPM_q_ivl_11886,
      b => LPM_q_ivl_11897,
      c => LPM_d0_ivl_11905
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3546
  U3414: xor_HPC2
    port map (
      a => LPM_q_ivl_11911,
      b => LPM_q_ivl_11922,
      c => LPM_d0_ivl_11930
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3547
  U3415: xnor_HPC2
    port map (
      a => LPM_q_ivl_11938,
      b => LPM_q_ivl_11945,
      c => LPM_d0_ivl_11953
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3548
  U3416: xnor_HPC2
    port map (
      a => LPM_q_ivl_11957,
      b => LPM_q_ivl_11964,
      c => LPM_d0_ivl_11972
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3549
  U3417: xnor_HPC2
    port map (
      a => LPM_q_ivl_11976,
      b => LPM_q_ivl_11983,
      c => LPM_d0_ivl_11991
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3550
  U3418: xor_HPC2
    port map (
      a => LPM_q_ivl_11997,
      b => LPM_q_ivl_12008,
      c => LPM_d0_ivl_12016
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3551
  U3419: xor_HPC2
    port map (
      a => LPM_q_ivl_12022,
      b => LPM_q_ivl_12029,
      c => LPM_d0_ivl_12037
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3072
  U3420: xnor_HPC2
    port map (
      a => LPM_q_ivl_3827,
      b => LPM_q_ivl_3838,
      c => LPM_d0_ivl_3846
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3552
  U3421: xnor_HPC2
    port map (
      a => LPM_q_ivl_12041,
      b => LPM_q_ivl_12048,
      c => LPM_d0_ivl_12056
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3553
  U3422: xnor_HPC2
    port map (
      a => LPM_q_ivl_12060,
      b => LPM_q_ivl_12067,
      c => LPM_d0_ivl_12079
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3554
  U3423: xnor_HPC2
    port map (
      a => LPM_q_ivl_12083,
      b => LPM_q_ivl_12090,
      c => LPM_d0_ivl_12098
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3555
  U3424: xnor_HPC2
    port map (
      a => LPM_q_ivl_12106,
      b => LPM_q_ivl_12115,
      c => LPM_d0_ivl_12123
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3556
  U3425: xnor_HPC2
    port map (
      a => LPM_q_ivl_12131,
      b => LPM_q_ivl_12138,
      c => LPM_d0_ivl_12146
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3557
  U3426: xnor_HPC2
    port map (
      a => LPM_q_ivl_12150,
      b => LPM_q_ivl_12157,
      c => LPM_d0_ivl_12169
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3558
  U3427: xor_HPC2
    port map (
      a => LPM_q_ivl_12175,
      b => LPM_q_ivl_12186,
      c => LPM_d0_ivl_12194
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3559
  U3428: xnor_HPC2
    port map (
      a => LPM_q_ivl_12198,
      b => LPM_q_ivl_12205,
      c => LPM_d0_ivl_12213
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3560
  U3429: xor_HPC2
    port map (
      a => LPM_q_ivl_12219,
      b => LPM_q_ivl_12230,
      c => LPM_d0_ivl_12238
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3561
  U3430: xnor_HPC2
    port map (
      a => LPM_q_ivl_12242,
      b => LPM_q_ivl_12249,
      c => LPM_d0_ivl_12257
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3562
  U3431: xnor_HPC2
    port map (
      a => LPM_q_ivl_12261,
      b => LPM_q_ivl_12268,
      c => LPM_d0_ivl_12276
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3563
  U3432: xnor_HPC2
    port map (
      a => LPM_q_ivl_12280,
      b => LPM_q_ivl_12287,
      c => LPM_d0_ivl_12295
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3564
  U3433: xnor_HPC2
    port map (
      a => LPM_q_ivl_12299,
      b => LPM_q_ivl_12306,
      c => LPM_d0_ivl_12318
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3565
  U3434: xnor_HPC2
    port map (
      a => LPM_q_ivl_12326,
      b => LPM_q_ivl_12335,
      c => LPM_d0_ivl_12343
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3566
  U3435: xnor_HPC2
    port map (
      a => LPM_q_ivl_12351,
      b => LPM_q_ivl_12358,
      c => LPM_d0_ivl_12366
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3567
  U3436: xnor_HPC2
    port map (
      a => LPM_q_ivl_12370,
      b => LPM_q_ivl_12377,
      c => LPM_d0_ivl_12385
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3568
  U3437: xnor_HPC2
    port map (
      a => LPM_q_ivl_12393,
      b => LPM_q_ivl_12402,
      c => LPM_d0_ivl_12410
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3569
  U3438: xnor_HPC2
    port map (
      a => LPM_q_ivl_12418,
      b => LPM_q_ivl_12425,
      c => LPM_d0_ivl_12433
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3570
  U3439: xnor_HPC2
    port map (
      a => LPM_q_ivl_12437,
      b => LPM_q_ivl_12444,
      c => LPM_d0_ivl_12456
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3571
  U3440: xnor_HPC2
    port map (
      a => LPM_q_ivl_12460,
      b => LPM_q_ivl_12467,
      c => LPM_d0_ivl_12475
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3572
  U3441: xnor_HPC2
    port map (
      a => LPM_q_ivl_12479,
      b => LPM_q_ivl_12486,
      c => LPM_d0_ivl_12498
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3573
  U3442: xnor_HPC2
    port map (
      a => LPM_q_ivl_12502,
      b => LPM_q_ivl_12509,
      c => LPM_d0_ivl_12517
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3574
  U3443: xnor_HPC2
    port map (
      a => LPM_q_ivl_12525,
      b => LPM_q_ivl_12534,
      c => LPM_d0_ivl_12542
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3575
  U3444: xnor_HPC2
    port map (
      a => LPM_q_ivl_12550,
      b => LPM_q_ivl_12557,
      c => LPM_d0_ivl_12565
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3576
  U3445: xnor_HPC2
    port map (
      a => LPM_q_ivl_12569,
      b => LPM_q_ivl_12576,
      c => LPM_d0_ivl_12588
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3577
  U3446: xor_HPC2
    port map (
      a => LPM_q_ivl_12594,
      b => LPM_q_ivl_12605,
      c => LPM_d0_ivl_12613
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3578
  U3447: xor_HPC2
    port map (
      a => LPM_q_ivl_12619,
      b => LPM_q_ivl_12630,
      c => LPM_d0_ivl_12638
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3579
  U3448: xnor_HPC2
    port map (
      a => LPM_q_ivl_12646,
      b => LPM_q_ivl_12653,
      c => LPM_d0_ivl_12661
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3580
  U3449: xnor_HPC2
    port map (
      a => LPM_q_ivl_12665,
      b => LPM_q_ivl_12672,
      c => LPM_d0_ivl_12680
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3581
  U3450: xnor_HPC2
    port map (
      a => LPM_q_ivl_12684,
      b => LPM_q_ivl_12691,
      c => LPM_d0_ivl_12699
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3582
  U3451: xor_HPC2
    port map (
      a => LPM_q_ivl_12705,
      b => LPM_q_ivl_12716,
      c => LPM_d0_ivl_12724
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3583
  U3452: xor_HPC2
    port map (
      a => LPM_q_ivl_12730,
      b => LPM_q_ivl_12741,
      c => LPM_d0_ivl_12749
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3584
  U3453: xnor_HPC2
    port map (
      a => LPM_q_ivl_12757,
      b => LPM_q_ivl_12764,
      c => LPM_d0_ivl_12772
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3585
  U3454: xnor_HPC2
    port map (
      a => LPM_q_ivl_12776,
      b => LPM_q_ivl_12783,
      c => LPM_d0_ivl_12791
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3586
  U3455: xnor_HPC2
    port map (
      a => LPM_q_ivl_12795,
      b => LPM_q_ivl_12802,
      c => LPM_d0_ivl_12814
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3587
  U3456: xor_HPC2
    port map (
      a => LPM_q_ivl_12820,
      b => LPM_q_ivl_12831,
      c => LPM_d0_ivl_12839
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3588
  U3457: xor_HPC2
    port map (
      a => LPM_q_ivl_12845,
      b => LPM_q_ivl_12852,
      c => LPM_d0_ivl_12860
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3073
  U3458: xnor_HPC2
    port map (
      a => LPM_q_ivl_3854,
      b => LPM_q_ivl_3865,
      c => LPM_d0_ivl_3873
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3589
  U3459: xnor_HPC2
    port map (
      a => LPM_q_ivl_12864,
      b => LPM_q_ivl_12871,
      c => LPM_d0_ivl_12879
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3590
  U3460: xor_HPC2
    port map (
      a => LPM_q_ivl_12885,
      b => LPM_q_ivl_12892,
      c => LPM_d0_ivl_12900
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3074
  U3461: xnor_HPC2
    port map (
      a => LPM_q_ivl_3881,
      b => LPM_q_ivl_3892,
      c => LPM_d0_ivl_3900
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3591
  U3462: xnor_HPC2
    port map (
      a => LPM_q_ivl_12904,
      b => LPM_q_ivl_12911,
      c => LPM_d0_ivl_12919
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3592
  U3463: xnor_HPC2
    port map (
      a => LPM_q_ivl_12923,
      b => LPM_q_ivl_12930,
      c => LPM_d0_ivl_12938
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3593
  U3464: xor_HPC2
    port map (
      a => LPM_q_ivl_12944,
      b => LPM_q_ivl_12955,
      c => LPM_d0_ivl_12963
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3594
  U3465: xor_HPC2
    port map (
      a => LPM_q_ivl_12969,
      b => LPM_q_ivl_12980,
      c => LPM_d0_ivl_12988
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3595
  U3466: xnor_HPC2
    port map (
      a => LPM_q_ivl_12996,
      b => LPM_q_ivl_13003,
      c => LPM_d0_ivl_13011
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3596
  U3467: xnor_HPC2
    port map (
      a => LPM_q_ivl_13015,
      b => LPM_q_ivl_13022,
      c => LPM_d0_ivl_13030
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3597
  U3468: xnor_HPC2
    port map (
      a => LPM_q_ivl_13034,
      b => LPM_q_ivl_13041,
      c => LPM_d0_ivl_13053
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3598
  U3469: xnor_HPC2
    port map (
      a => LPM_q_ivl_13057,
      b => LPM_q_ivl_13064,
      c => LPM_d0_ivl_13072
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3599
  U3470: xnor_HPC2
    port map (
      a => LPM_q_ivl_13080,
      b => LPM_q_ivl_13089,
      c => LPM_d0_ivl_13097
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3600
  U3471: xnor_HPC2
    port map (
      a => LPM_q_ivl_13105,
      b => LPM_q_ivl_13112,
      c => LPM_d0_ivl_13120
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3601
  U3472: xnor_HPC2
    port map (
      a => LPM_q_ivl_13124,
      b => LPM_q_ivl_13131,
      c => LPM_d0_ivl_13143
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3602
  U3473: xnor_HPC2
    port map (
      a => LPM_q_ivl_13147,
      b => LPM_q_ivl_13154,
      c => LPM_d0_ivl_13162
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3603
  U3474: xnor_HPC2
    port map (
      a => LPM_q_ivl_13170,
      b => LPM_q_ivl_13179,
      c => LPM_d0_ivl_13187
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3604
  U3475: xnor_HPC2
    port map (
      a => LPM_q_ivl_13195,
      b => LPM_q_ivl_13202,
      c => LPM_d0_ivl_13210
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3605
  U3476: xnor_HPC2
    port map (
      a => LPM_q_ivl_13214,
      b => LPM_q_ivl_13221,
      c => LPM_d0_ivl_13233
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3606
  U3477: xnor_HPC2
    port map (
      a => LPM_q_ivl_13237,
      b => LPM_q_ivl_13244,
      c => LPM_d0_ivl_13252
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3607
  U3478: xnor_HPC2
    port map (
      a => LPM_q_ivl_13256,
      b => LPM_q_ivl_13263,
      c => LPM_d0_ivl_13275
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3608
  U3479: xor_HPC2
    port map (
      a => LPM_q_ivl_13281,
      b => LPM_q_ivl_13292,
      c => LPM_d0_ivl_13300
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3609
  U3480: xor_HPC2
    port map (
      a => LPM_q_ivl_13306,
      b => LPM_q_ivl_13317,
      c => LPM_d0_ivl_13325
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3610
  U3481: xnor_HPC2
    port map (
      a => LPM_q_ivl_13333,
      b => LPM_q_ivl_13340,
      c => LPM_d0_ivl_13348
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3611
  U3482: xnor_HPC2
    port map (
      a => LPM_q_ivl_13352,
      b => LPM_q_ivl_13359,
      c => LPM_d0_ivl_13367
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3612
  U3483: xnor_HPC2
    port map (
      a => LPM_q_ivl_13371,
      b => LPM_q_ivl_13378,
      c => LPM_d0_ivl_13386
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3613
  U3484: xor_HPC2
    port map (
      a => LPM_q_ivl_13392,
      b => LPM_q_ivl_13403,
      c => LPM_d0_ivl_13411
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3614
  U3485: xor_HPC2
    port map (
      a => LPM_q_ivl_13417,
      b => LPM_q_ivl_13428,
      c => LPM_d0_ivl_13436
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3615
  U3486: xnor_HPC2
    port map (
      a => LPM_q_ivl_13444,
      b => LPM_q_ivl_13451,
      c => LPM_d0_ivl_13459
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3616
  U3487: xnor_HPC2
    port map (
      a => LPM_q_ivl_13463,
      b => LPM_q_ivl_13470,
      c => LPM_d0_ivl_13478
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3617
  U3488: xnor_HPC2
    port map (
      a => LPM_q_ivl_13482,
      b => LPM_q_ivl_13489,
      c => LPM_d0_ivl_13501
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3618
  U3489: xor_HPC2
    port map (
      a => LPM_q_ivl_13507,
      b => LPM_q_ivl_13518,
      c => LPM_d0_ivl_13526
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3619
  U3490: xor_HPC2
    port map (
      a => LPM_q_ivl_13532,
      b => LPM_q_ivl_13543,
      c => LPM_d0_ivl_13551
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3620
  U3491: xnor_HPC2
    port map (
      a => LPM_q_ivl_13559,
      b => LPM_q_ivl_13566,
      c => LPM_d0_ivl_13574
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3621
  U3492: xnor_HPC2
    port map (
      a => LPM_q_ivl_13578,
      b => LPM_q_ivl_13585,
      c => LPM_d0_ivl_13593
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3622
  U3493: xor_HPC2
    port map (
      a => LPM_q_ivl_13599,
      b => LPM_q_ivl_13610,
      c => LPM_d0_ivl_13618
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3623
  U3494: xor_HPC2
    port map (
      a => LPM_q_ivl_13624,
      b => LPM_q_ivl_13631,
      c => LPM_d0_ivl_13639
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3075
  U3495: xnor_HPC2
    port map (
      a => LPM_q_ivl_3908,
      b => LPM_q_ivl_3919,
      c => LPM_d0_ivl_3927
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3624
  U3496: xnor_HPC2
    port map (
      a => LPM_q_ivl_13643,
      b => LPM_q_ivl_13650,
      c => LPM_d0_ivl_13658
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3625
  U3497: xnor_HPC2
    port map (
      a => LPM_q_ivl_13662,
      b => LPM_q_ivl_13669,
      c => LPM_d0_ivl_13677
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3626
  U3498: xor_HPC2
    port map (
      a => LPM_q_ivl_13683,
      b => LPM_q_ivl_13694,
      c => LPM_d0_ivl_13702
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3627
  U3499: xor_HPC2
    port map (
      a => LPM_q_ivl_13708,
      b => LPM_q_ivl_13715,
      c => LPM_d0_ivl_13723
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3076
  U3500: xnor_HPC2
    port map (
      a => LPM_q_ivl_3935,
      b => LPM_q_ivl_3946,
      c => LPM_d0_ivl_3954
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3628
  U3501: xnor_HPC2
    port map (
      a => LPM_q_ivl_13727,
      b => LPM_q_ivl_13734,
      c => LPM_d0_ivl_13742
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3629
  U3502: xnor_HPC2
    port map (
      a => LPM_q_ivl_13746,
      b => LPM_q_ivl_13753,
      c => LPM_d0_ivl_13765
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3630
  U3503: xnor_HPC2
    port map (
      a => LPM_q_ivl_13769,
      b => LPM_q_ivl_13776,
      c => LPM_d0_ivl_13784
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3631
  U3504: xnor_HPC2
    port map (
      a => LPM_q_ivl_13792,
      b => LPM_q_ivl_13801,
      c => LPM_d0_ivl_13809
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3632
  U3505: xnor_HPC2
    port map (
      a => LPM_q_ivl_13817,
      b => LPM_q_ivl_13824,
      c => LPM_d0_ivl_13832
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3633
  U3506: xnor_HPC2
    port map (
      a => LPM_q_ivl_13836,
      b => LPM_q_ivl_13843,
      c => LPM_d0_ivl_13855
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3634
  U3507: xnor_HPC2
    port map (
      a => LPM_q_ivl_13859,
      b => LPM_q_ivl_13866,
      c => LPM_d0_ivl_13874
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3635
  U3508: xnor_HPC2
    port map (
      a => LPM_q_ivl_13878,
      b => LPM_q_ivl_13885,
      c => LPM_d0_ivl_13897
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3636
  U3509: xnor_HPC2
    port map (
      a => LPM_q_ivl_13901,
      b => LPM_q_ivl_13908,
      c => LPM_d0_ivl_13916
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3637
  U3510: xnor_HPC2
    port map (
      a => LPM_q_ivl_13920,
      b => LPM_q_ivl_13927,
      c => LPM_d0_ivl_13935
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3638
  U3511: xor_HPC2
    port map (
      a => LPM_q_ivl_13941,
      b => LPM_q_ivl_13952,
      c => LPM_d0_ivl_13960
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3639
  U3512: xnor_HPC2
    port map (
      a => LPM_q_ivl_13964,
      b => LPM_q_ivl_13971,
      c => LPM_d0_ivl_13979
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3640
  U3513: xnor_HPC2
    port map (
      a => LPM_q_ivl_13983,
      b => LPM_q_ivl_13990,
      c => LPM_d0_ivl_14002
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3641
  U3514: xor_HPC2
    port map (
      a => LPM_q_ivl_14008,
      b => LPM_q_ivl_14019,
      c => LPM_d0_ivl_14027
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3642
  U3515: xnor_HPC2
    port map (
      a => LPM_q_ivl_14035,
      b => LPM_q_ivl_14042,
      c => LPM_d0_ivl_14050
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3643
  U3516: xnor_HPC2
    port map (
      a => LPM_q_ivl_14054,
      b => LPM_q_ivl_14061,
      c => LPM_d0_ivl_14069
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3644
  U3517: xnor_HPC2
    port map (
      a => LPM_q_ivl_14073,
      b => LPM_q_ivl_14080,
      c => LPM_d0_ivl_14088
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3645
  U3518: xor_HPC2
    port map (
      a => LPM_q_ivl_14094,
      b => LPM_q_ivl_14105,
      c => LPM_d0_ivl_14113
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3646
  U3519: xor_HPC2
    port map (
      a => LPM_q_ivl_14119,
      b => LPM_q_ivl_14130,
      c => LPM_d0_ivl_14138
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3647
  U3520: xnor_HPC2
    port map (
      a => LPM_q_ivl_14146,
      b => LPM_q_ivl_14153,
      c => LPM_d0_ivl_14161
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3648
  U3521: xnor_HPC2
    port map (
      a => LPM_q_ivl_14165,
      b => LPM_q_ivl_14172,
      c => LPM_d0_ivl_14180
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3649
  U3522: xnor_HPC2
    port map (
      a => LPM_q_ivl_14184,
      b => LPM_q_ivl_14191,
      c => LPM_d0_ivl_14203
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3650
  U3523: xor_HPC2
    port map (
      a => LPM_q_ivl_14209,
      b => LPM_q_ivl_14220,
      c => LPM_d0_ivl_14228
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3651
  U3524: xnor_HPC2
    port map (
      a => LPM_q_ivl_14232,
      b => LPM_q_ivl_14239,
      c => LPM_d0_ivl_14247
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3652
  U3525: xor_HPC2
    port map (
      a => LPM_q_ivl_14253,
      b => LPM_q_ivl_14264,
      c => LPM_d0_ivl_14272
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3653
  U3526: xnor_HPC2
    port map (
      a => LPM_q_ivl_14276,
      b => LPM_q_ivl_14283,
      c => LPM_d0_ivl_14291
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3654
  U3527: xnor_HPC2
    port map (
      a => LPM_q_ivl_14295,
      b => LPM_q_ivl_14302,
      c => LPM_d0_ivl_14310
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3655
  U3528: xnor_HPC2
    port map (
      a => LPM_q_ivl_14314,
      b => LPM_q_ivl_14321,
      c => LPM_d0_ivl_14329
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3656
  U3529: xnor_HPC2
    port map (
      a => LPM_q_ivl_14333,
      b => LPM_q_ivl_14340,
      c => LPM_d0_ivl_14352
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3657
  U3530: xor_HPC2
    port map (
      a => LPM_q_ivl_14358,
      b => LPM_q_ivl_14369,
      c => LPM_d0_ivl_14377
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3658
  U3531: xnor_HPC2
    port map (
      a => LPM_q_ivl_14385,
      b => LPM_q_ivl_14392,
      c => LPM_d0_ivl_14400
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3659
  U3532: xnor_HPC2
    port map (
      a => LPM_q_ivl_14404,
      b => LPM_q_ivl_14411,
      c => LPM_d0_ivl_14419
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3660
  U3533: xnor_HPC2
    port map (
      a => LPM_q_ivl_14423,
      b => LPM_q_ivl_14430,
      c => LPM_d0_ivl_14438
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3661
  U3534: xor_HPC2
    port map (
      a => LPM_q_ivl_14444,
      b => LPM_q_ivl_14455,
      c => LPM_d0_ivl_14463
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3662
  U3535: xnor_HPC2
    port map (
      a => LPM_q_ivl_14471,
      b => LPM_q_ivl_14478,
      c => LPM_d0_ivl_14486
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3663
  U3536: xnor_HPC2
    port map (
      a => LPM_q_ivl_14490,
      b => LPM_q_ivl_14497,
      c => LPM_d0_ivl_14505
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3664
  U3537: xnor_HPC2
    port map (
      a => LPM_q_ivl_14509,
      b => LPM_q_ivl_14516,
      c => LPM_d0_ivl_14528
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3665
  U3538: xnor_HPC2
    port map (
      a => LPM_q_ivl_14532,
      b => LPM_q_ivl_14539,
      c => LPM_d0_ivl_14547
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3666
  U3539: xnor_HPC2
    port map (
      a => LPM_q_ivl_14551,
      b => LPM_q_ivl_14558,
      c => LPM_d0_ivl_14570
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3667
  U3540: xor_HPC2
    port map (
      a => LPM_q_ivl_14576,
      b => LPM_q_ivl_14587,
      c => LPM_d0_ivl_14595
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3668
  U3541: xnor_HPC2
    port map (
      a => LPM_q_ivl_14603,
      b => LPM_q_ivl_14612,
      c => LPM_d0_ivl_14620
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3669
  U3542: xnor_HPC2
    port map (
      a => LPM_q_ivl_14624,
      b => LPM_q_ivl_14631,
      c => LPM_d0_ivl_14639
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3670
  U3543: xor_HPC2
    port map (
      a => LPM_q_ivl_14645,
      b => LPM_q_ivl_14656,
      c => LPM_d0_ivl_14664
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3671
  U3544: xnor_HPC2
    port map (
      a => LPM_q_ivl_14668,
      b => LPM_q_ivl_14675,
      c => LPM_d0_ivl_14683
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3672
  U3545: xnor_HPC2
    port map (
      a => LPM_q_ivl_14687,
      b => LPM_q_ivl_14694,
      c => LPM_d0_ivl_14702
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3673
  U3546: xnor_HPC2
    port map (
      a => LPM_q_ivl_14706,
      b => LPM_q_ivl_14713,
      c => LPM_d0_ivl_14721
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3674
  U3547: xnor_HPC2
    port map (
      a => LPM_q_ivl_14725,
      b => LPM_q_ivl_14732,
      c => LPM_d0_ivl_14744
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3675
  U3548: xnor_HPC2
    port map (
      a => LPM_q_ivl_14748,
      b => LPM_q_ivl_14755,
      c => LPM_d0_ivl_14763
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3676
  U3549: xnor_HPC2
    port map (
      a => LPM_q_ivl_14771,
      b => LPM_q_ivl_14778,
      c => LPM_d0_ivl_14786
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3677
  U3550: xnor_HPC2
    port map (
      a => LPM_q_ivl_14790,
      b => LPM_q_ivl_14797,
      c => LPM_d0_ivl_14809
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3678
  U3551: xor_HPC2
    port map (
      a => LPM_q_ivl_14815,
      b => LPM_q_ivl_14826,
      c => LPM_d0_ivl_14834
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3679
  U3552: xor_HPC2
    port map (
      a => LPM_q_ivl_14840,
      b => LPM_q_ivl_14851,
      c => LPM_d0_ivl_14859
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3680
  U3553: xnor_HPC2
    port map (
      a => LPM_q_ivl_14867,
      b => LPM_q_ivl_14874,
      c => LPM_d0_ivl_14882
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3681
  U3554: xnor_HPC2
    port map (
      a => LPM_q_ivl_14886,
      b => LPM_q_ivl_14893,
      c => LPM_d0_ivl_14901
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3682
  U3555: xor_HPC2
    port map (
      a => LPM_q_ivl_14907,
      b => LPM_q_ivl_14918,
      c => LPM_d0_ivl_14926
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3683
  U3556: xnor_HPC2
    port map (
      a => LPM_q_ivl_14934,
      b => LPM_q_ivl_14941,
      c => LPM_d0_ivl_14949
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3684
  U3557: xnor_HPC2
    port map (
      a => LPM_q_ivl_14953,
      b => LPM_q_ivl_14960,
      c => LPM_d0_ivl_14968
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3685
  U3558: xnor_HPC2
    port map (
      a => LPM_q_ivl_14972,
      b => LPM_q_ivl_14979,
      c => LPM_d0_ivl_14987
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3686
  U3559: xor_HPC2
    port map (
      a => LPM_q_ivl_14993,
      b => LPM_q_ivl_15004,
      c => LPM_d0_ivl_15012
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3687
  U3560: xor_HPC2
    port map (
      a => LPM_q_ivl_15018,
      b => LPM_q_ivl_15025,
      c => LPM_d0_ivl_15033
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3077
  U3561: xnor_HPC2
    port map (
      a => LPM_q_ivl_3962,
      b => LPM_q_ivl_3973,
      c => LPM_d0_ivl_3981
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3688
  U3562: xnor_HPC2
    port map (
      a => LPM_q_ivl_15037,
      b => LPM_q_ivl_15044,
      c => LPM_d0_ivl_15052
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3689
  U3563: xnor_HPC2
    port map (
      a => LPM_q_ivl_15056,
      b => LPM_q_ivl_15063,
      c => LPM_d0_ivl_15075
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3690
  U3564: xnor_HPC2
    port map (
      a => LPM_q_ivl_15079,
      b => LPM_q_ivl_15086,
      c => LPM_d0_ivl_15094
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3691
  U3565: xnor_HPC2
    port map (
      a => LPM_q_ivl_15098,
      b => LPM_q_ivl_15105,
      c => LPM_d0_ivl_15117
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3692
  U3566: xnor_HPC2
    port map (
      a => LPM_q_ivl_15121,
      b => LPM_q_ivl_15128,
      c => LPM_d0_ivl_15136
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3693
  U3567: xnor_HPC2
    port map (
      a => LPM_q_ivl_15140,
      b => LPM_q_ivl_15147,
      c => LPM_d0_ivl_15159
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3694
  U3568: xor_HPC2
    port map (
      a => LPM_q_ivl_15165,
      b => LPM_q_ivl_15176,
      c => LPM_d0_ivl_15184
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3695
  U3569: xnor_HPC2
    port map (
      a => LPM_q_ivl_15188,
      b => LPM_q_ivl_15195,
      c => LPM_d0_ivl_15203
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3696
  U3570: xnor_HPC2
    port map (
      a => LPM_q_ivl_15207,
      b => LPM_q_ivl_15214,
      c => LPM_d0_ivl_15222
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3697
  U3571: xnor_HPC2
    port map (
      a => LPM_q_ivl_15226,
      b => LPM_q_ivl_15233,
      c => LPM_d0_ivl_15241
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3698
  U3572: xnor_HPC2
    port map (
      a => LPM_q_ivl_15245,
      b => LPM_q_ivl_15252,
      c => LPM_d0_ivl_15260
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3699
  U3573: xnor_HPC2
    port map (
      a => LPM_q_ivl_15264,
      b => LPM_q_ivl_15271,
      c => LPM_d0_ivl_15283
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3700
  U3574: xor_HPC2
    port map (
      a => LPM_q_ivl_15289,
      b => LPM_q_ivl_15300,
      c => LPM_d0_ivl_15308
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3701
  U3575: xnor_HPC2
    port map (
      a => LPM_q_ivl_15316,
      b => LPM_q_ivl_15323,
      c => LPM_d0_ivl_15331
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3702
  U3576: xnor_HPC2
    port map (
      a => LPM_q_ivl_15335,
      b => LPM_q_ivl_15342,
      c => LPM_d0_ivl_15350
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3703
  U3577: xnor_HPC2
    port map (
      a => LPM_q_ivl_15354,
      b => LPM_q_ivl_15361,
      c => LPM_d0_ivl_15369
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3704
  U3578: xor_HPC2
    port map (
      a => LPM_q_ivl_15375,
      b => LPM_q_ivl_15382,
      c => LPM_d0_ivl_15390
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3078
  U3579: xnor_HPC2
    port map (
      a => LPM_q_ivl_3989,
      b => LPM_q_ivl_4000,
      c => LPM_d0_ivl_4008
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3705
  U3580: xnor_HPC2
    port map (
      a => LPM_q_ivl_15394,
      b => LPM_q_ivl_15401,
      c => LPM_d0_ivl_15409
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3706
  U3581: xnor_HPC2
    port map (
      a => LPM_q_ivl_15413,
      b => LPM_q_ivl_15420,
      c => LPM_d0_ivl_15432
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3707
  U3582: xnor_HPC2
    port map (
      a => LPM_q_ivl_15436,
      b => LPM_q_ivl_15443,
      c => LPM_d0_ivl_15451
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3708
  U3583: xnor_HPC2
    port map (
      a => LPM_q_ivl_15455,
      b => LPM_q_ivl_15462,
      c => LPM_d0_ivl_15474
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3709
  U3584: xnor_HPC2
    port map (
      a => LPM_q_ivl_15478,
      b => LPM_q_ivl_15485,
      c => LPM_d0_ivl_15493
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3710
  U3585: xnor_HPC2
    port map (
      a => LPM_q_ivl_15501,
      b => LPM_q_ivl_15510,
      c => LPM_d0_ivl_15518
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3711
  U3586: xnor_HPC2
    port map (
      a => LPM_q_ivl_15526,
      b => LPM_q_ivl_15533,
      c => LPM_d0_ivl_15541
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3712
  U3587: xnor_HPC2
    port map (
      a => LPM_q_ivl_15545,
      b => LPM_q_ivl_15552,
      c => LPM_d0_ivl_15564
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3713
  U3588: xnor_HPC2
    port map (
      a => LPM_q_ivl_15568,
      b => LPM_q_ivl_15575,
      c => LPM_d0_ivl_15583
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3714
  U3589: xnor_HPC2
    port map (
      a => LPM_q_ivl_15587,
      b => LPM_q_ivl_15594,
      c => LPM_d0_ivl_15606
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3715
  U3590: xnor_HPC2
    port map (
      a => LPM_q_ivl_15610,
      b => LPM_q_ivl_15617,
      c => LPM_d0_ivl_15625
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3716
  U3591: xnor_HPC2
    port map (
      a => LPM_q_ivl_15629,
      b => LPM_q_ivl_15636,
      c => LPM_d0_ivl_15648
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3717
  U3592: xnor_HPC2
    port map (
      a => LPM_q_ivl_15652,
      b => LPM_q_ivl_15659,
      c => LPM_d0_ivl_15667
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3718
  U3593: xor_HPC2
    port map (
      a => LPM_q_ivl_15673,
      b => LPM_q_ivl_15684,
      c => LPM_d0_ivl_15692
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3719
  U3594: xor_HPC2
    port map (
      a => LPM_q_ivl_15698,
      b => LPM_q_ivl_15709,
      c => LPM_d0_ivl_15717
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3720
  U3595: xnor_HPC2
    port map (
      a => LPM_q_ivl_15725,
      b => LPM_q_ivl_15732,
      c => LPM_d0_ivl_15740
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3721
  U3596: xnor_HPC2
    port map (
      a => LPM_q_ivl_15744,
      b => LPM_q_ivl_15751,
      c => LPM_d0_ivl_15759
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3722
  U3597: xnor_HPC2
    port map (
      a => LPM_q_ivl_15763,
      b => LPM_q_ivl_15770,
      c => LPM_d0_ivl_15782
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3723
  U3598: xnor_HPC2
    port map (
      a => LPM_q_ivl_15786,
      b => LPM_q_ivl_15793,
      c => LPM_d0_ivl_15801
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3724
  U3599: xor_HPC2
    port map (
      a => LPM_q_ivl_15807,
      b => LPM_q_ivl_15818,
      c => LPM_d0_ivl_15826
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3725
  U3600: xor_HPC2
    port map (
      a => LPM_q_ivl_15832,
      b => LPM_q_ivl_15843,
      c => LPM_d0_ivl_15851
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3726
  U3601: xnor_HPC2
    port map (
      a => LPM_q_ivl_15859,
      b => LPM_q_ivl_15866,
      c => LPM_d0_ivl_15874
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3727
  U3602: xnor_HPC2
    port map (
      a => LPM_q_ivl_15878,
      b => LPM_q_ivl_15885,
      c => LPM_d0_ivl_15893
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3728
  U3603: xnor_HPC2
    port map (
      a => LPM_q_ivl_15897,
      b => LPM_q_ivl_15904,
      c => LPM_d0_ivl_15916
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3729
  U3604: xnor_HPC2
    port map (
      a => LPM_q_ivl_15920,
      b => LPM_q_ivl_15927,
      c => LPM_d0_ivl_15935
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3730
  U3605: xor_HPC2
    port map (
      a => LPM_q_ivl_15941,
      b => LPM_q_ivl_15952,
      c => LPM_d0_ivl_15960
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3731
  U3606: xor_HPC2
    port map (
      a => LPM_q_ivl_15966,
      b => LPM_q_ivl_15973,
      c => LPM_d0_ivl_15981
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3079
  U3607: xnor_HPC2
    port map (
      a => LPM_q_ivl_4016,
      b => LPM_q_ivl_4027,
      c => LPM_d0_ivl_4035
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3732
  U3608: xnor_HPC2
    port map (
      a => LPM_q_ivl_15985,
      b => LPM_q_ivl_15992,
      c => LPM_d0_ivl_16000
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3733
  U3609: xnor_HPC2
    port map (
      a => LPM_q_ivl_16004,
      b => LPM_q_ivl_16011,
      c => LPM_d0_ivl_16023
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3734
  U3610: xnor_HPC2
    port map (
      a => LPM_q_ivl_16027,
      b => LPM_q_ivl_16034,
      c => LPM_d0_ivl_16042
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3735
  U3611: xnor_HPC2
    port map (
      a => LPM_q_ivl_16046,
      b => LPM_q_ivl_16053,
      c => LPM_d0_ivl_16065
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3736
  U3612: xnor_HPC2
    port map (
      a => LPM_q_ivl_16069,
      b => LPM_q_ivl_16076,
      c => LPM_d0_ivl_16084
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3737
  U3613: xnor_HPC2
    port map (
      a => LPM_q_ivl_16092,
      b => LPM_q_ivl_16101,
      c => LPM_d0_ivl_16109
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3738
  U3614: xnor_HPC2
    port map (
      a => LPM_q_ivl_16113,
      b => LPM_q_ivl_16120,
      c => LPM_d0_ivl_16128
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3739
  U3615: xnor_HPC2
    port map (
      a => LPM_q_ivl_16132,
      b => LPM_q_ivl_16139,
      c => LPM_d0_ivl_16151
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3740
  U3616: xor_HPC2
    port map (
      a => LPM_q_ivl_16157,
      b => LPM_q_ivl_16168,
      c => LPM_d0_ivl_16176
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3741
  U3617: xnor_HPC2
    port map (
      a => LPM_q_ivl_16180,
      b => LPM_q_ivl_16187,
      c => LPM_d0_ivl_16195
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3742
  U3618: xnor_HPC2
    port map (
      a => LPM_q_ivl_16199,
      b => LPM_q_ivl_16206,
      c => LPM_d0_ivl_16214
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3743
  U3619: xnor_HPC2
    port map (
      a => LPM_q_ivl_16218,
      b => LPM_q_ivl_16225,
      c => LPM_d0_ivl_16233
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3744
  U3620: xnor_HPC2
    port map (
      a => LPM_q_ivl_16237,
      b => LPM_q_ivl_16244,
      c => LPM_d0_ivl_16256
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3745
  U3621: xnor_HPC2
    port map (
      a => LPM_q_ivl_16260,
      b => LPM_q_ivl_16267,
      c => LPM_d0_ivl_16275
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3746
  U3622: xnor_HPC2
    port map (
      a => LPM_q_ivl_16283,
      b => LPM_q_ivl_16290,
      c => LPM_d0_ivl_16298
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3747
  U3623: xnor_HPC2
    port map (
      a => LPM_q_ivl_16302,
      b => LPM_q_ivl_16309,
      c => LPM_d0_ivl_16321
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3748
  U3624: xor_HPC2
    port map (
      a => LPM_q_ivl_16327,
      b => LPM_q_ivl_16338,
      c => LPM_d0_ivl_16346
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3749
  U3625: xnor_HPC2
    port map (
      a => LPM_q_ivl_16350,
      b => LPM_q_ivl_16357,
      c => LPM_d0_ivl_16365
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3750
  U3626: xnor_HPC2
    port map (
      a => LPM_q_ivl_16369,
      b => LPM_q_ivl_16376,
      c => LPM_d0_ivl_16384
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3751
  U3627: xnor_HPC2
    port map (
      a => LPM_q_ivl_16388,
      b => LPM_q_ivl_16395,
      c => LPM_d0_ivl_16403
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3752
  U3628: xor_HPC2
    port map (
      a => LPM_q_ivl_16409,
      b => LPM_q_ivl_16420,
      c => LPM_d0_ivl_16428
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3753
  U3629: xnor_HPC2
    port map (
      a => LPM_q_ivl_16432,
      b => LPM_q_ivl_16439,
      c => LPM_d0_ivl_16447
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3754
  U3630: xnor_HPC2
    port map (
      a => LPM_q_ivl_16451,
      b => LPM_q_ivl_16458,
      c => LPM_d0_ivl_16470
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3755
  U3631: xnor_HPC2
    port map (
      a => LPM_q_ivl_16474,
      b => LPM_q_ivl_16481,
      c => LPM_d0_ivl_16489
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3756
  U3632: xor_HPC2
    port map (
      a => LPM_q_ivl_16495,
      b => LPM_q_ivl_16506,
      c => LPM_d0_ivl_16514
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3757
  U3633: xnor_HPC2
    port map (
      a => LPM_q_ivl_16522,
      b => LPM_q_ivl_16529,
      c => LPM_d0_ivl_16537
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3758
  U3634: xnor_HPC2
    port map (
      a => LPM_q_ivl_16541,
      b => LPM_q_ivl_16548,
      c => LPM_d0_ivl_16556
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3759
  U3635: xnor_HPC2
    port map (
      a => LPM_q_ivl_16560,
      b => LPM_q_ivl_16567,
      c => LPM_d0_ivl_16579
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3760
  U3636: xor_HPC2
    port map (
      a => LPM_q_ivl_16585,
      b => LPM_q_ivl_16596,
      c => LPM_d0_ivl_16604
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3761
  U3637: xnor_HPC2
    port map (
      a => LPM_q_ivl_16608,
      b => LPM_q_ivl_16615,
      c => LPM_d0_ivl_16623
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3762
  U3638: xnor_HPC2
    port map (
      a => LPM_q_ivl_16627,
      b => LPM_q_ivl_16634,
      c => LPM_d0_ivl_16642
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3763
  U3639: xnor_HPC2
    port map (
      a => LPM_q_ivl_16646,
      b => LPM_q_ivl_16653,
      c => LPM_d0_ivl_16661
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3764
  U3640: xnor_HPC2
    port map (
      a => LPM_q_ivl_16665,
      b => LPM_q_ivl_16672,
      c => LPM_d0_ivl_16680
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3765
  U3641: xnor_HPC2
    port map (
      a => LPM_q_ivl_16684,
      b => LPM_q_ivl_16691,
      c => LPM_d0_ivl_16703
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3766
  U3642: xor_HPC2
    port map (
      a => LPM_q_ivl_16709,
      b => LPM_q_ivl_16720,
      c => LPM_d0_ivl_16728
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3767
  U3643: xnor_HPC2
    port map (
      a => LPM_q_ivl_16736,
      b => LPM_q_ivl_16743,
      c => LPM_d0_ivl_16751
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3768
  U3644: xnor_HPC2
    port map (
      a => LPM_q_ivl_16755,
      b => LPM_q_ivl_16762,
      c => LPM_d0_ivl_16770
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3769
  U3645: xnor_HPC2
    port map (
      a => LPM_q_ivl_16774,
      b => LPM_q_ivl_16781,
      c => LPM_d0_ivl_16789
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3770
  U3646: xor_HPC2
    port map (
      a => LPM_q_ivl_16795,
      b => LPM_q_ivl_16806,
      c => LPM_d0_ivl_16814
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3771
  U3647: xnor_HPC2
    port map (
      a => LPM_q_ivl_16822,
      b => LPM_q_ivl_16829,
      c => LPM_d0_ivl_16837
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3772
  U3648: xnor_HPC2
    port map (
      a => LPM_q_ivl_16841,
      b => LPM_q_ivl_16848,
      c => LPM_d0_ivl_16856
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3773
  U3649: xnor_HPC2
    port map (
      a => LPM_q_ivl_16860,
      b => LPM_q_ivl_16867,
      c => LPM_d0_ivl_16879
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3774
  U3650: xnor_HPC2
    port map (
      a => LPM_q_ivl_16883,
      b => LPM_q_ivl_16890,
      c => LPM_d0_ivl_16898
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3775
  U3651: xnor_HPC2
    port map (
      a => LPM_q_ivl_16902,
      b => LPM_q_ivl_16909,
      c => LPM_d0_ivl_16921
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3776
  U3652: xnor_HPC2
    port map (
      a => LPM_q_ivl_16925,
      b => LPM_q_ivl_16932,
      c => LPM_d0_ivl_16940
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3777
  U3653: xnor_HPC2
    port map (
      a => LPM_q_ivl_16948,
      b => LPM_q_ivl_16957,
      c => LPM_d0_ivl_16965
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3778
  U3654: xnor_HPC2
    port map (
      a => LPM_q_ivl_16973,
      b => LPM_q_ivl_16980,
      c => LPM_d0_ivl_16988
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3779
  U3655: xnor_HPC2
    port map (
      a => LPM_q_ivl_16992,
      b => LPM_q_ivl_16999,
      c => LPM_d0_ivl_17011
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3780
  U3656: xnor_HPC2
    port map (
      a => LPM_q_ivl_17015,
      b => LPM_q_ivl_17022,
      c => LPM_d0_ivl_17030
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3781
  U3657: xnor_HPC2
    port map (
      a => LPM_q_ivl_17034,
      b => LPM_q_ivl_17041,
      c => LPM_d0_ivl_17053
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3782
  U3658: xnor_HPC2
    port map (
      a => LPM_q_ivl_17057,
      b => LPM_q_ivl_17064,
      c => LPM_d0_ivl_17072
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3783
  U3659: xnor_HPC2
    port map (
      a => LPM_q_ivl_17076,
      b => LPM_q_ivl_17083,
      c => LPM_d0_ivl_17095
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3784
  U3660: xnor_HPC2
    port map (
      a => LPM_q_ivl_17099,
      b => LPM_q_ivl_17106,
      c => LPM_d0_ivl_17114
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3785
  U3661: xor_HPC2
    port map (
      a => LPM_q_ivl_17120,
      b => LPM_q_ivl_17131,
      c => LPM_d0_ivl_17139
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3786
  U3662: xor_HPC2
    port map (
      a => LPM_q_ivl_17145,
      b => LPM_q_ivl_17156,
      c => LPM_d0_ivl_17164
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3787
  U3663: xnor_HPC2
    port map (
      a => LPM_q_ivl_17172,
      b => LPM_q_ivl_17179,
      c => LPM_d0_ivl_17187
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3788
  U3664: xnor_HPC2
    port map (
      a => LPM_q_ivl_17191,
      b => LPM_q_ivl_17198,
      c => LPM_d0_ivl_17206
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3789
  U3665: xnor_HPC2
    port map (
      a => LPM_q_ivl_17210,
      b => LPM_q_ivl_17217,
      c => LPM_d0_ivl_17229
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3790
  U3666: xnor_HPC2
    port map (
      a => LPM_q_ivl_17233,
      b => LPM_q_ivl_17240,
      c => LPM_d0_ivl_17248
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3791
  U3667: xor_HPC2
    port map (
      a => LPM_q_ivl_17254,
      b => LPM_q_ivl_17265,
      c => LPM_d0_ivl_17273
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3792
  U3668: xor_HPC2
    port map (
      a => LPM_q_ivl_17279,
      b => LPM_q_ivl_17286,
      c => LPM_d0_ivl_17294
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3080
  U3669: xnor_HPC2
    port map (
      a => LPM_q_ivl_4043,
      b => LPM_q_ivl_4054,
      c => LPM_d0_ivl_4062
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3793
  U3670: xnor_HPC2
    port map (
      a => LPM_q_ivl_17298,
      b => LPM_q_ivl_17305,
      c => LPM_d0_ivl_17313
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3794
  U3671: xnor_HPC2
    port map (
      a => LPM_q_ivl_17317,
      b => LPM_q_ivl_17324,
      c => LPM_d0_ivl_17336
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3795
  U3672: xnor_HPC2
    port map (
      a => LPM_q_ivl_17340,
      b => LPM_q_ivl_17347,
      c => LPM_d0_ivl_17355
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3796
  U3673: xnor_HPC2
    port map (
      a => LPM_q_ivl_17359,
      b => LPM_q_ivl_17366,
      c => LPM_d0_ivl_17378
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3797
  U3674: xor_HPC2
    port map (
      a => LPM_q_ivl_17384,
      b => LPM_q_ivl_17395,
      c => LPM_d0_ivl_17403
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3798
  U3675: xnor_HPC2
    port map (
      a => LPM_q_ivl_17407,
      b => LPM_q_ivl_17414,
      c => LPM_d0_ivl_17422
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3799
  U3676: xnor_HPC2
    port map (
      a => LPM_q_ivl_17426,
      b => LPM_q_ivl_17433,
      c => LPM_d0_ivl_17441
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3800
  U3677: xnor_HPC2
    port map (
      a => LPM_q_ivl_17445,
      b => LPM_q_ivl_17452,
      c => LPM_d0_ivl_17460
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3801
  U3678: xnor_HPC2
    port map (
      a => LPM_q_ivl_17464,
      b => LPM_q_ivl_17471,
      c => LPM_d0_ivl_17483
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3802
  U3679: xnor_HPC2
    port map (
      a => LPM_q_ivl_17487,
      b => LPM_q_ivl_17494,
      c => LPM_d0_ivl_17502
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3803
  U3680: xor_HPC2
    port map (
      a => LPM_q_ivl_17508,
      b => LPM_q_ivl_17519,
      c => LPM_d0_ivl_17527
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3804
  U3681: xnor_HPC2
    port map (
      a => LPM_q_ivl_17535,
      b => LPM_q_ivl_17542,
      c => LPM_d0_ivl_17550
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3805
  U3682: xnor_HPC2
    port map (
      a => LPM_q_ivl_17554,
      b => LPM_q_ivl_17561,
      c => LPM_d0_ivl_17569
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3806
  U3683: xnor_HPC2
    port map (
      a => LPM_q_ivl_17573,
      b => LPM_q_ivl_17580,
      c => LPM_d0_ivl_17592
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3807
  U3684: xnor_HPC2
    port map (
      a => LPM_q_ivl_17596,
      b => LPM_q_ivl_17603,
      c => LPM_d0_ivl_17611
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3808
  U3685: xnor_HPC2
    port map (
      a => LPM_q_ivl_17619,
      b => LPM_q_ivl_17628,
      c => LPM_d0_ivl_17636
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3809
  U3686: xnor_HPC2
    port map (
      a => LPM_q_ivl_17640,
      b => LPM_q_ivl_17647,
      c => LPM_d0_ivl_17655
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3810
  U3687: xnor_HPC2
    port map (
      a => LPM_q_ivl_17659,
      b => LPM_q_ivl_17666,
      c => LPM_d0_ivl_17678
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3811
  U3688: xnor_HPC2
    port map (
      a => LPM_q_ivl_17682,
      b => LPM_q_ivl_17689,
      c => LPM_d0_ivl_17697
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3812
  U3689: xnor_HPC2
    port map (
      a => LPM_q_ivl_17701,
      b => LPM_q_ivl_17708,
      c => LPM_d0_ivl_17720
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3813
  U3690: xnor_HPC2
    port map (
      a => LPM_q_ivl_17724,
      b => LPM_q_ivl_17731,
      c => LPM_d0_ivl_17739
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3814
  U3691: xnor_HPC2
    port map (
      a => LPM_q_ivl_17747,
      b => LPM_q_ivl_17754,
      c => LPM_d0_ivl_17762
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3815
  U3692: xnor_HPC2
    port map (
      a => LPM_q_ivl_17766,
      b => LPM_q_ivl_17773,
      c => LPM_d0_ivl_17785
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3816
  U3693: xnor_HPC2
    port map (
      a => LPM_q_ivl_17789,
      b => LPM_q_ivl_17796,
      c => LPM_d0_ivl_17804
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3817
  U3694: xor_HPC2
    port map (
      a => LPM_q_ivl_17810,
      b => LPM_q_ivl_17821,
      c => LPM_d0_ivl_17829
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3818
  U3695: xor_HPC2
    port map (
      a => LPM_q_ivl_17835,
      b => LPM_q_ivl_17846,
      c => LPM_d0_ivl_17854
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3819
  U3696: xnor_HPC2
    port map (
      a => LPM_q_ivl_17862,
      b => LPM_q_ivl_17869,
      c => LPM_d0_ivl_17877
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3820
  U3697: xnor_HPC2
    port map (
      a => LPM_q_ivl_17881,
      b => LPM_q_ivl_17888,
      c => LPM_d0_ivl_17896
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3821
  U3698: xnor_HPC2
    port map (
      a => LPM_q_ivl_17900,
      b => LPM_q_ivl_17907,
      c => LPM_d0_ivl_17919
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3822
  U3699: xnor_HPC2
    port map (
      a => LPM_q_ivl_17923,
      b => LPM_q_ivl_17930,
      c => LPM_d0_ivl_17938
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3823
  U3700: xor_HPC2
    port map (
      a => LPM_q_ivl_17944,
      b => LPM_q_ivl_17951,
      c => LPM_d0_ivl_17959
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3081
  U3701: xnor_HPC2
    port map (
      a => LPM_q_ivl_4070,
      b => LPM_q_ivl_4081,
      c => LPM_d0_ivl_4089
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3824
  U3702: xnor_HPC2
    port map (
      a => LPM_q_ivl_17963,
      b => LPM_q_ivl_17970,
      c => LPM_d0_ivl_17978
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3825
  U3703: xnor_HPC2
    port map (
      a => LPM_q_ivl_17982,
      b => LPM_q_ivl_17989,
      c => LPM_d0_ivl_18001
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3826
  U3704: xor_HPC2
    port map (
      a => LPM_q_ivl_18007,
      b => LPM_q_ivl_18018,
      c => LPM_d0_ivl_18026
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3827
  U3705: xnor_HPC2
    port map (
      a => LPM_q_ivl_18030,
      b => LPM_q_ivl_18037,
      c => LPM_d0_ivl_18045
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3828
  U3706: xnor_HPC2
    port map (
      a => LPM_q_ivl_18049,
      b => LPM_q_ivl_18056,
      c => LPM_d0_ivl_18064
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3829
  U3707: xnor_HPC2
    port map (
      a => LPM_q_ivl_18068,
      b => LPM_q_ivl_18075,
      c => LPM_d0_ivl_18083
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3830
  U3708: xnor_HPC2
    port map (
      a => LPM_q_ivl_18087,
      b => LPM_q_ivl_18094,
      c => LPM_d0_ivl_18106
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3831
  U3709: xnor_HPC2
    port map (
      a => LPM_q_ivl_18110,
      b => LPM_q_ivl_18117,
      c => LPM_d0_ivl_18125
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3832
  U3710: xor_HPC2
    port map (
      a => LPM_q_ivl_18131,
      b => LPM_q_ivl_18142,
      c => LPM_d0_ivl_18150
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3833
  U3711: xnor_HPC2
    port map (
      a => LPM_q_ivl_18158,
      b => LPM_q_ivl_18165,
      c => LPM_d0_ivl_18173
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3834
  U3712: xnor_HPC2
    port map (
      a => LPM_q_ivl_18177,
      b => LPM_q_ivl_18184,
      c => LPM_d0_ivl_18192
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3835
  U3713: xnor_HPC2
    port map (
      a => LPM_q_ivl_18196,
      b => LPM_q_ivl_18203,
      c => LPM_d0_ivl_18215
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3836
  U3714: xnor_HPC2
    port map (
      a => LPM_q_ivl_18219,
      b => LPM_q_ivl_18226,
      c => LPM_d0_ivl_18234
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3837
  U3715: xnor_HPC2
    port map (
      a => LPM_q_ivl_18242,
      b => LPM_q_ivl_18251,
      c => LPM_d0_ivl_18259
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3838
  U3716: xnor_HPC2
    port map (
      a => LPM_q_ivl_18267,
      b => LPM_q_ivl_18274,
      c => LPM_d0_ivl_18282
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3839
  U3717: xnor_HPC2
    port map (
      a => LPM_q_ivl_18286,
      b => LPM_q_ivl_18293,
      c => LPM_d0_ivl_18305
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3840
  U3718: xnor_HPC2
    port map (
      a => LPM_q_ivl_18309,
      b => LPM_q_ivl_18316,
      c => LPM_d0_ivl_18324
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3841
  U3719: xnor_HPC2
    port map (
      a => LPM_q_ivl_18328,
      b => LPM_q_ivl_18335,
      c => LPM_d0_ivl_18347
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3842
  U3720: xnor_HPC2
    port map (
      a => LPM_q_ivl_18351,
      b => LPM_q_ivl_18358,
      c => LPM_d0_ivl_18366
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3843
  U3721: xnor_HPC2
    port map (
      a => LPM_q_ivl_18370,
      b => LPM_q_ivl_18377,
      c => LPM_d0_ivl_18389
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3844
  U3722: xor_HPC2
    port map (
      a => LPM_q_ivl_18395,
      b => LPM_q_ivl_18406,
      c => LPM_d0_ivl_18414
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3845
  U3723: xnor_HPC2
    port map (
      a => LPM_q_ivl_18418,
      b => LPM_q_ivl_18425,
      c => LPM_d0_ivl_18433
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3846
  U3724: xnor_HPC2
    port map (
      a => LPM_q_ivl_18437,
      b => LPM_q_ivl_18444,
      c => LPM_d0_ivl_18452
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3847
  U3725: xnor_HPC2
    port map (
      a => LPM_q_ivl_18456,
      b => LPM_q_ivl_18463,
      c => LPM_d0_ivl_18471
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3848
  U3726: xnor_HPC2
    port map (
      a => LPM_q_ivl_18475,
      b => LPM_q_ivl_18482,
      c => LPM_d0_ivl_18490
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3849
  U3727: xnor_HPC2
    port map (
      a => LPM_q_ivl_18494,
      b => LPM_q_ivl_18501,
      c => LPM_d0_ivl_18513
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3850
  U3728: xnor_HPC2
    port map (
      a => LPM_q_ivl_18517,
      b => LPM_q_ivl_18524,
      c => LPM_d0_ivl_18532
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3851
  U3729: xor_HPC2
    port map (
      a => LPM_q_ivl_18538,
      b => LPM_q_ivl_18549,
      c => LPM_d0_ivl_18557
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3852
  U3730: xnor_HPC2
    port map (
      a => LPM_q_ivl_18565,
      b => LPM_q_ivl_18572,
      c => LPM_d0_ivl_18580
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3853
  U3731: xnor_HPC2
    port map (
      a => LPM_q_ivl_18584,
      b => LPM_q_ivl_18591,
      c => LPM_d0_ivl_18599
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3854
  U3732: xnor_HPC2
    port map (
      a => LPM_q_ivl_18603,
      b => LPM_q_ivl_18610,
      c => LPM_d0_ivl_18622
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3855
  U3733: xnor_HPC2
    port map (
      a => LPM_q_ivl_18626,
      b => LPM_q_ivl_18633,
      c => LPM_d0_ivl_18641
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3856
  U3734: xor_HPC2
    port map (
      a => LPM_q_ivl_18647,
      b => LPM_q_ivl_18658,
      c => LPM_d0_ivl_18666
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3857
  U3735: xor_HPC2
    port map (
      a => LPM_q_ivl_18672,
      b => LPM_q_ivl_18683,
      c => LPM_d0_ivl_18691
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3858
  U3736: xnor_HPC2
    port map (
      a => LPM_q_ivl_18699,
      b => LPM_q_ivl_18706,
      c => LPM_d0_ivl_18714
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3859
  U3737: xnor_HPC2
    port map (
      a => LPM_q_ivl_18718,
      b => LPM_q_ivl_18725,
      c => LPM_d0_ivl_18733
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3860
  U3738: xnor_HPC2
    port map (
      a => LPM_q_ivl_18737,
      b => LPM_q_ivl_18744,
      c => LPM_d0_ivl_18756
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3861
  U3739: xnor_HPC2
    port map (
      a => LPM_q_ivl_18760,
      b => LPM_q_ivl_18767,
      c => LPM_d0_ivl_18775
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3862
  U3740: xnor_HPC2
    port map (
      a => LPM_q_ivl_18779,
      b => LPM_q_ivl_18786,
      c => LPM_d0_ivl_18794
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3863
  U3741: xnor_HPC2
    port map (
      a => LPM_q_ivl_18798,
      b => LPM_q_ivl_18805,
      c => LPM_d0_ivl_18813
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3864
  U3742: xor_HPC2
    port map (
      a => LPM_q_ivl_18819,
      b => LPM_q_ivl_18830,
      c => LPM_d0_ivl_18838
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3865
  U3743: xnor_HPC2
    port map (
      a => LPM_q_ivl_18842,
      b => LPM_q_ivl_18849,
      c => LPM_d0_ivl_18857
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3866
  U3744: xnor_HPC2
    port map (
      a => LPM_q_ivl_18861,
      b => LPM_q_ivl_18868,
      c => LPM_d0_ivl_18880
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3867
  U3745: xnor_HPC2
    port map (
      a => LPM_q_ivl_18884,
      b => LPM_q_ivl_18891,
      c => LPM_d0_ivl_18899
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3868
  U3746: xor_HPC2
    port map (
      a => LPM_q_ivl_18905,
      b => LPM_q_ivl_18916,
      c => LPM_d0_ivl_18924
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3869
  U3747: xnor_HPC2
    port map (
      a => LPM_q_ivl_18932,
      b => LPM_q_ivl_18939,
      c => LPM_d0_ivl_18947
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3870
  U3748: xnor_HPC2
    port map (
      a => LPM_q_ivl_18951,
      b => LPM_q_ivl_18958,
      c => LPM_d0_ivl_18966
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3871
  U3749: xnor_HPC2
    port map (
      a => LPM_q_ivl_18970,
      b => LPM_q_ivl_18977,
      c => LPM_d0_ivl_18989
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3872
  U3750: xnor_HPC2
    port map (
      a => LPM_q_ivl_18993,
      b => LPM_q_ivl_19000,
      c => LPM_d0_ivl_19008
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3873
  U3751: xor_HPC2
    port map (
      a => LPM_q_ivl_19014,
      b => LPM_q_ivl_19025,
      c => LPM_d0_ivl_19033
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3874
  U3752: xnor_HPC2
    port map (
      a => LPM_q_ivl_19041,
      b => LPM_q_ivl_19048,
      c => LPM_d0_ivl_19056
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3875
  U3753: xnor_HPC2
    port map (
      a => LPM_q_ivl_19060,
      b => LPM_q_ivl_19067,
      c => LPM_d0_ivl_19075
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3876
  U3754: xnor_HPC2
    port map (
      a => LPM_q_ivl_19079,
      b => LPM_q_ivl_19086,
      c => LPM_d0_ivl_19098
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3877
  U3755: xnor_HPC2
    port map (
      a => LPM_q_ivl_19106,
      b => LPM_q_ivl_19115,
      c => LPM_d0_ivl_19123
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3878
  U3756: xnor_HPC2
    port map (
      a => LPM_q_ivl_19127,
      b => LPM_q_ivl_19134,
      c => LPM_d0_ivl_19142
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3879
  U3757: xnor_HPC2
    port map (
      a => LPM_q_ivl_19146,
      b => LPM_q_ivl_19153,
      c => LPM_d0_ivl_19161
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3880
  U3758: xnor_HPC2
    port map (
      a => LPM_q_ivl_19165,
      b => LPM_q_ivl_19172,
      c => LPM_d0_ivl_19180
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3881
  U3759: xnor_HPC2
    port map (
      a => LPM_q_ivl_19184,
      b => LPM_q_ivl_19191,
      c => LPM_d0_ivl_19199
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3882
  U3760: xnor_HPC2
    port map (
      a => LPM_q_ivl_19203,
      b => LPM_q_ivl_19210,
      c => LPM_d0_ivl_19222
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3883
  U3761: xnor_HPC2
    port map (
      a => LPM_q_ivl_19226,
      b => LPM_q_ivl_19233,
      c => LPM_d0_ivl_19241
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3884
  U3762: xnor_HPC2
    port map (
      a => LPM_q_ivl_19249,
      b => LPM_q_ivl_19256,
      c => LPM_d0_ivl_19264
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3885
  U3763: xnor_HPC2
    port map (
      a => LPM_q_ivl_19268,
      b => LPM_q_ivl_19275,
      c => LPM_d0_ivl_19287
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3886
  U3764: xnor_HPC2
    port map (
      a => LPM_q_ivl_19291,
      b => LPM_q_ivl_19298,
      c => LPM_d0_ivl_19306
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3887
  U3765: xnor_HPC2
    port map (
      a => LPM_q_ivl_19310,
      b => LPM_q_ivl_19317,
      c => LPM_d0_ivl_19325
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3888
  U3766: xor_HPC2
    port map (
      a => LPM_q_ivl_19331,
      b => LPM_q_ivl_19342,
      c => LPM_d0_ivl_19350
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3889
  U3767: xnor_HPC2
    port map (
      a => LPM_q_ivl_19354,
      b => LPM_q_ivl_19361,
      c => LPM_d0_ivl_19369
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3890
  U3768: xnor_HPC2
    port map (
      a => LPM_q_ivl_19373,
      b => LPM_q_ivl_19380,
      c => LPM_d0_ivl_19392
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3891
  U3769: xnor_HPC2
    port map (
      a => LPM_q_ivl_19396,
      b => LPM_q_ivl_19403,
      c => LPM_d0_ivl_19411
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3892
  U3770: xor_HPC2
    port map (
      a => LPM_q_ivl_19417,
      b => LPM_q_ivl_19424,
      c => LPM_d0_ivl_19432
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3082
  U3771: xnor_HPC2
    port map (
      a => LPM_q_ivl_4097,
      b => LPM_q_ivl_4108,
      c => LPM_d0_ivl_4116
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3893
  U3772: xnor_HPC2
    port map (
      a => LPM_q_ivl_19436,
      b => LPM_q_ivl_19443,
      c => LPM_d0_ivl_19451
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3894
  U3773: xnor_HPC2
    port map (
      a => LPM_q_ivl_19455,
      b => LPM_q_ivl_19462,
      c => LPM_d0_ivl_19474
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3895
  U3774: xnor_HPC2
    port map (
      a => LPM_q_ivl_19478,
      b => LPM_q_ivl_19485,
      c => LPM_d0_ivl_19493
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3896
  U3775: xnor_HPC2
    port map (
      a => LPM_q_ivl_19497,
      b => LPM_q_ivl_19504,
      c => LPM_d0_ivl_19512
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3897
  U3776: xor_HPC2
    port map (
      a => LPM_q_ivl_19518,
      b => LPM_q_ivl_19529,
      c => LPM_d0_ivl_19537
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3898
  U3777: xnor_HPC2
    port map (
      a => LPM_q_ivl_19541,
      b => LPM_q_ivl_19548,
      c => LPM_d0_ivl_19556
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3899
  U3778: xnor_HPC2
    port map (
      a => LPM_q_ivl_19560,
      b => LPM_q_ivl_19567,
      c => LPM_d0_ivl_19579
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3900
  U3779: xnor_HPC2
    port map (
      a => LPM_q_ivl_19583,
      b => LPM_q_ivl_19590,
      c => LPM_d0_ivl_19598
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3901
  U3780: xor_HPC2
    port map (
      a => LPM_q_ivl_19604,
      b => LPM_q_ivl_19615,
      c => LPM_d0_ivl_19623
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3902
  U3781: xnor_HPC2
    port map (
      a => LPM_q_ivl_19631,
      b => LPM_q_ivl_19638,
      c => LPM_d0_ivl_19646
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3903
  U3782: xnor_HPC2
    port map (
      a => LPM_q_ivl_19650,
      b => LPM_q_ivl_19657,
      c => LPM_d0_ivl_19665
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3904
  U3783: xnor_HPC2
    port map (
      a => LPM_q_ivl_19669,
      b => LPM_q_ivl_19676,
      c => LPM_d0_ivl_19688
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3905
  U3784: xnor_HPC2
    port map (
      a => LPM_q_ivl_19692,
      b => LPM_q_ivl_19699,
      c => LPM_d0_ivl_19707
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3906
  U3785: xnor_HPC2
    port map (
      a => LPM_q_ivl_19715,
      b => LPM_q_ivl_19724,
      c => LPM_d0_ivl_19732
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3907
  U3786: xnor_HPC2
    port map (
      a => LPM_q_ivl_19736,
      b => LPM_q_ivl_19743,
      c => LPM_d0_ivl_19751
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3908
  U3787: xnor_HPC2
    port map (
      a => LPM_q_ivl_19755,
      b => LPM_q_ivl_19762,
      c => LPM_d0_ivl_19774
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3909
  U3788: xnor_HPC2
    port map (
      a => LPM_q_ivl_19778,
      b => LPM_q_ivl_19785,
      c => LPM_d0_ivl_19793
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3910
  U3789: xnor_HPC2
    port map (
      a => LPM_q_ivl_19801,
      b => LPM_q_ivl_19808,
      c => LPM_d0_ivl_19816
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3911
  U3790: xnor_HPC2
    port map (
      a => LPM_q_ivl_19820,
      b => LPM_q_ivl_19827,
      c => LPM_d0_ivl_19839
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3912
  U3791: xnor_HPC2
    port map (
      a => LPM_q_ivl_19843,
      b => LPM_q_ivl_19850,
      c => LPM_d0_ivl_19858
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3913
  U3792: xnor_HPC2
    port map (
      a => LPM_q_ivl_19862,
      b => LPM_q_ivl_19869,
      c => LPM_d0_ivl_19881
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3914
  U3793: xnor_HPC2
    port map (
      a => LPM_q_ivl_19885,
      b => LPM_q_ivl_19892,
      c => LPM_d0_ivl_19900
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3915
  U3794: xnor_HPC2
    port map (
      a => LPM_q_ivl_19904,
      b => LPM_q_ivl_19911,
      c => LPM_d0_ivl_19923
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3916
  U3795: xnor_HPC2
    port map (
      a => LPM_q_ivl_19927,
      b => LPM_q_ivl_19934,
      c => LPM_d0_ivl_19942
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3917
  U3796: xor_HPC2
    port map (
      a => LPM_q_ivl_19948,
      b => LPM_q_ivl_19959,
      c => LPM_d0_ivl_19967
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3918
  U3797: xnor_HPC2
    port map (
      a => LPM_q_ivl_19971,
      b => LPM_q_ivl_19978,
      c => LPM_d0_ivl_19986
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3919
  U3798: xnor_HPC2
    port map (
      a => LPM_q_ivl_19990,
      b => LPM_q_ivl_19997,
      c => LPM_d0_ivl_20009
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3920
  U3799: xnor_HPC2
    port map (
      a => LPM_q_ivl_20013,
      b => LPM_q_ivl_20020,
      c => LPM_d0_ivl_20028
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3921
  U3800: xnor_HPC2
    port map (
      a => LPM_q_ivl_20032,
      b => LPM_q_ivl_20039,
      c => LPM_d0_ivl_20051
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3922
  U3801: xnor_HPC2
    port map (
      a => LPM_q_ivl_20055,
      b => LPM_q_ivl_20062,
      c => LPM_d0_ivl_20070
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3923
  U3802: xor_HPC2
    port map (
      a => LPM_q_ivl_20076,
      b => LPM_q_ivl_20087,
      c => LPM_d0_ivl_20095
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3924
  U3803: xnor_HPC2
    port map (
      a => LPM_q_ivl_20103,
      b => LPM_q_ivl_20110,
      c => LPM_d0_ivl_20118
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3925
  U3804: xnor_HPC2
    port map (
      a => LPM_q_ivl_20122,
      b => LPM_q_ivl_20129,
      c => LPM_d0_ivl_20137
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3926
  U3805: xnor_HPC2
    port map (
      a => LPM_q_ivl_20141,
      b => LPM_q_ivl_20148,
      c => LPM_d0_ivl_20160
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3927
  U3806: xnor_HPC2
    port map (
      a => LPM_q_ivl_20164,
      b => LPM_q_ivl_20171,
      c => LPM_d0_ivl_20179
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3928
  U3807: xnor_HPC2
    port map (
      a => LPM_q_ivl_20183,
      b => LPM_q_ivl_20190,
      c => LPM_d0_ivl_20202
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3929
  U3808: xnor_HPC2
    port map (
      a => LPM_q_ivl_20206,
      b => LPM_q_ivl_20213,
      c => LPM_d0_ivl_20221
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3930
  U3809: xor_HPC2
    port map (
      a => LPM_q_ivl_20227,
      b => LPM_q_ivl_20238,
      c => LPM_d0_ivl_20246
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3931
  U3810: xnor_HPC2
    port map (
      a => LPM_q_ivl_20250,
      b => LPM_q_ivl_20257,
      c => LPM_d0_ivl_20265
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3932
  U3811: xnor_HPC2
    port map (
      a => LPM_q_ivl_20269,
      b => LPM_q_ivl_20276,
      c => LPM_d0_ivl_20288
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3933
  U3812: xnor_HPC2
    port map (
      a => LPM_q_ivl_20292,
      b => LPM_q_ivl_20299,
      c => LPM_d0_ivl_20307
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3934
  U3813: xor_HPC2
    port map (
      a => LPM_q_ivl_20313,
      b => LPM_q_ivl_20324,
      c => LPM_d0_ivl_20332
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3935
  U3814: xnor_HPC2
    port map (
      a => LPM_q_ivl_20340,
      b => LPM_q_ivl_20347,
      c => LPM_d0_ivl_20355
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3936
  U3815: xnor_HPC2
    port map (
      a => LPM_q_ivl_20359,
      b => LPM_q_ivl_20366,
      c => LPM_d0_ivl_20374
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3937
  U3816: xnor_HPC2
    port map (
      a => LPM_q_ivl_20378,
      b => LPM_q_ivl_20385,
      c => LPM_d0_ivl_20397
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3938
  U3817: xnor_HPC2
    port map (
      a => LPM_q_ivl_20401,
      b => LPM_q_ivl_20408,
      c => LPM_d0_ivl_20416
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3939
  U3818: xnor_HPC2
    port map (
      a => LPM_q_ivl_20424,
      b => LPM_q_ivl_20433,
      c => LPM_d0_ivl_20441
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3940
  U3819: xnor_HPC2
    port map (
      a => LPM_q_ivl_20445,
      b => LPM_q_ivl_20452,
      c => LPM_d0_ivl_20460
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3941
  U3820: xnor_HPC2
    port map (
      a => LPM_q_ivl_20464,
      b => LPM_q_ivl_20471,
      c => LPM_d0_ivl_20483
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3942
  U3821: xnor_HPC2
    port map (
      a => LPM_q_ivl_20487,
      b => LPM_q_ivl_20494,
      c => LPM_d0_ivl_20502
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3943
  U3822: xnor_HPC2
    port map (
      a => LPM_q_ivl_20506,
      b => LPM_q_ivl_20513,
      c => LPM_d0_ivl_20525
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3944
  U3823: xnor_HPC2
    port map (
      a => LPM_q_ivl_20529,
      b => LPM_q_ivl_20536,
      c => LPM_d0_ivl_20544
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3945
  U3824: xnor_HPC2
    port map (
      a => LPM_q_ivl_20552,
      b => LPM_q_ivl_20559,
      c => LPM_d0_ivl_20567
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3946
  U3825: xnor_HPC2
    port map (
      a => LPM_q_ivl_20571,
      b => LPM_q_ivl_20578,
      c => LPM_d0_ivl_20590
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3947
  U3826: xnor_HPC2
    port map (
      a => LPM_q_ivl_20594,
      b => LPM_q_ivl_20601,
      c => LPM_d0_ivl_20609
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3948
  U3827: xnor_HPC2
    port map (
      a => LPM_q_ivl_20613,
      b => LPM_q_ivl_20620,
      c => LPM_d0_ivl_20632
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3949
  U3828: xnor_HPC2
    port map (
      a => LPM_q_ivl_20636,
      b => LPM_q_ivl_20643,
      c => LPM_d0_ivl_20651
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3950
  U3829: xnor_HPC2
    port map (
      a => LPM_q_ivl_20655,
      b => LPM_q_ivl_20662,
      c => LPM_d0_ivl_20674
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3951
  U3830: xnor_HPC2
    port map (
      a => LPM_q_ivl_20678,
      b => LPM_q_ivl_20685,
      c => LPM_d0_ivl_20693
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3952
  U3831: xor_HPC2
    port map (
      a => LPM_q_ivl_20699,
      b => LPM_q_ivl_20710,
      c => LPM_d0_ivl_20718
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3953
  U3832: xnor_HPC2
    port map (
      a => LPM_q_ivl_20722,
      b => LPM_q_ivl_20729,
      c => LPM_d0_ivl_20737
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3954
  U3833: xnor_HPC2
    port map (
      a => LPM_q_ivl_20741,
      b => LPM_q_ivl_20748,
      c => LPM_d0_ivl_20760
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3955
  U3834: xnor_HPC2
    port map (
      a => LPM_q_ivl_20764,
      b => LPM_q_ivl_20771,
      c => LPM_d0_ivl_20779
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3956
  U3835: xnor_HPC2
    port map (
      a => LPM_q_ivl_20783,
      b => LPM_q_ivl_20790,
      c => LPM_d0_ivl_20802
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3957
  U3836: xnor_HPC2
    port map (
      a => LPM_q_ivl_20806,
      b => LPM_q_ivl_20813,
      c => LPM_d0_ivl_20821
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3958
  U3837: xor_HPC2
    port map (
      a => LPM_q_ivl_20827,
      b => LPM_q_ivl_20838,
      c => LPM_d0_ivl_20846
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3959
  U3838: xnor_HPC2
    port map (
      a => LPM_q_ivl_20854,
      b => LPM_q_ivl_20861,
      c => LPM_d0_ivl_20869
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3960
  U3839: xnor_HPC2
    port map (
      a => LPM_q_ivl_20873,
      b => LPM_q_ivl_20880,
      c => LPM_d0_ivl_20888
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3961
  U3840: xnor_HPC2
    port map (
      a => LPM_q_ivl_20892,
      b => LPM_q_ivl_20899,
      c => LPM_d0_ivl_20911
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3962
  U3841: xnor_HPC2
    port map (
      a => LPM_q_ivl_20915,
      b => LPM_q_ivl_20922,
      c => LPM_d0_ivl_20930
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3963
  U3842: xnor_HPC2
    port map (
      a => LPM_q_ivl_20934,
      b => LPM_q_ivl_20941,
      c => LPM_d0_ivl_20953
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3964
  U3843: xnor_HPC2
    port map (
      a => LPM_q_ivl_20957,
      b => LPM_q_ivl_20964,
      c => LPM_d0_ivl_20972
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3965
  U3844: xnor_HPC2
    port map (
      a => LPM_q_ivl_20980,
      b => LPM_q_ivl_20989,
      c => LPM_d0_ivl_20997
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3966
  U3845: xnor_HPC2
    port map (
      a => LPM_q_ivl_21001,
      b => LPM_q_ivl_21008,
      c => LPM_d0_ivl_21016
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3967
  U3846: xnor_HPC2
    port map (
      a => LPM_q_ivl_21020,
      b => LPM_q_ivl_21027,
      c => LPM_d0_ivl_21035
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3968
  U3847: xnor_HPC2
    port map (
      a => LPM_q_ivl_21039,
      b => LPM_q_ivl_21046,
      c => LPM_d0_ivl_21054
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3969
  U3848: xnor_HPC2
    port map (
      a => LPM_q_ivl_21058,
      b => LPM_q_ivl_21065,
      c => LPM_d0_ivl_21077
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3970
  U3849: xnor_HPC2
    port map (
      a => LPM_q_ivl_21081,
      b => LPM_q_ivl_21088,
      c => LPM_d0_ivl_21096
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3971
  U3850: xnor_HPC2
    port map (
      a => LPM_q_ivl_21104,
      b => LPM_q_ivl_21111,
      c => LPM_d0_ivl_21119
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3972
  U3851: xnor_HPC2
    port map (
      a => LPM_q_ivl_21123,
      b => LPM_q_ivl_21130,
      c => LPM_d0_ivl_21142
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3973
  U3852: xnor_HPC2
    port map (
      a => LPM_q_ivl_21146,
      b => LPM_q_ivl_21153,
      c => LPM_d0_ivl_21161
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3974
  U3853: xnor_HPC2
    port map (
      a => LPM_q_ivl_21165,
      b => LPM_q_ivl_21172,
      c => LPM_d0_ivl_21184
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3975
  U3854: xnor_HPC2
    port map (
      a => LPM_q_ivl_21188,
      b => LPM_q_ivl_21195,
      c => LPM_d0_ivl_21203
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3976
  U3855: xor_HPC2
    port map (
      a => LPM_q_ivl_21209,
      b => LPM_q_ivl_21220,
      c => LPM_d0_ivl_21228
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3977
  U3856: xnor_HPC2
    port map (
      a => LPM_q_ivl_21232,
      b => LPM_q_ivl_21239,
      c => LPM_d0_ivl_21247
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3978
  U3857: xnor_HPC2
    port map (
      a => LPM_q_ivl_21251,
      b => LPM_q_ivl_21258,
      c => LPM_d0_ivl_21270
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3979
  U3858: xnor_HPC2
    port map (
      a => LPM_q_ivl_21274,
      b => LPM_q_ivl_21281,
      c => LPM_d0_ivl_21289
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3980
  U3859: xnor_HPC2
    port map (
      a => LPM_q_ivl_21293,
      b => LPM_q_ivl_21300,
      c => LPM_d0_ivl_21312
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3981
  U3860: xnor_HPC2
    port map (
      a => LPM_q_ivl_21316,
      b => LPM_q_ivl_21323,
      c => LPM_d0_ivl_21331
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3982
  U3861: xnor_HPC2
    port map (
      a => LPM_q_ivl_21335,
      b => LPM_q_ivl_21342,
      c => LPM_d0_ivl_21354
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3983
  U3862: xnor_HPC2
    port map (
      a => LPM_q_ivl_21358,
      b => LPM_q_ivl_21365,
      c => LPM_d0_ivl_21373
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3984
  U3863: xor_HPC2
    port map (
      a => LPM_q_ivl_21379,
      b => LPM_q_ivl_21386,
      c => LPM_d0_ivl_21394
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3083
  U3864: xnor_HPC2
    port map (
      a => LPM_q_ivl_4124,
      b => LPM_q_ivl_4135,
      c => LPM_d0_ivl_4143
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3985
  U3865: xnor_HPC2
    port map (
      a => LPM_q_ivl_21398,
      b => LPM_q_ivl_21405,
      c => LPM_d0_ivl_21413
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3986
  U3866: xnor_HPC2
    port map (
      a => LPM_q_ivl_21417,
      b => LPM_q_ivl_21424,
      c => LPM_d0_ivl_21436
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3987
  U3867: xnor_HPC2
    port map (
      a => LPM_q_ivl_21440,
      b => LPM_q_ivl_21447,
      c => LPM_d0_ivl_21455
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3988
  U3868: xnor_HPC2
    port map (
      a => LPM_q_ivl_21459,
      b => LPM_q_ivl_21466,
      c => LPM_d0_ivl_21478
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3989
  U3869: xnor_HPC2
    port map (
      a => LPM_q_ivl_21482,
      b => LPM_q_ivl_21489,
      c => LPM_d0_ivl_21497
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3990
  U3870: xor_HPC2
    port map (
      a => LPM_q_ivl_21503,
      b => LPM_q_ivl_21514,
      c => LPM_d0_ivl_21522
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3991
  U3871: xnor_HPC2
    port map (
      a => LPM_q_ivl_21526,
      b => LPM_q_ivl_21533,
      c => LPM_d0_ivl_21541
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3992
  U3872: xnor_HPC2
    port map (
      a => LPM_q_ivl_21545,
      b => LPM_q_ivl_21552,
      c => LPM_d0_ivl_21564
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3993
  U3873: xnor_HPC2
    port map (
      a => LPM_q_ivl_21568,
      b => LPM_q_ivl_21575,
      c => LPM_d0_ivl_21583
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3994
  U3874: xnor_HPC2
    port map (
      a => LPM_q_ivl_21587,
      b => LPM_q_ivl_21594,
      c => LPM_d0_ivl_21606
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3995
  U3875: xnor_HPC2
    port map (
      a => LPM_q_ivl_21610,
      b => LPM_q_ivl_21617,
      c => LPM_d0_ivl_21625
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3996
  U3876: xnor_HPC2
    port map (
      a => LPM_q_ivl_21629,
      b => LPM_q_ivl_21636,
      c => LPM_d0_ivl_21648
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3997
  U3877: xnor_HPC2
    port map (
      a => LPM_q_ivl_21652,
      b => LPM_q_ivl_21659,
      c => LPM_d0_ivl_21667
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3998
  U3878: xor_HPC2
    port map (
      a => LPM_q_ivl_21673,
      b => LPM_q_ivl_21684,
      c => LPM_d0_ivl_21692
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3999
  U3879: xnor_HPC2
    port map (
      a => LPM_q_ivl_21700,
      b => LPM_q_ivl_21707,
      c => LPM_d0_ivl_21715
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4000
  U3880: xnor_HPC2
    port map (
      a => LPM_q_ivl_21719,
      b => LPM_q_ivl_21726,
      c => LPM_d0_ivl_21734
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4001
  U3881: xnor_HPC2
    port map (
      a => LPM_q_ivl_21738,
      b => LPM_q_ivl_21745,
      c => LPM_d0_ivl_21757
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4002
  U3882: xnor_HPC2
    port map (
      a => LPM_q_ivl_21761,
      b => LPM_q_ivl_21768,
      c => LPM_d0_ivl_21776
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4003
  U3883: xnor_HPC2
    port map (
      a => LPM_q_ivl_21780,
      b => LPM_q_ivl_21787,
      c => LPM_d0_ivl_21799
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4004
  U3884: xnor_HPC2
    port map (
      a => LPM_q_ivl_21803,
      b => LPM_q_ivl_21810,
      c => LPM_d0_ivl_21818
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4005
  U3885: xnor_HPC2
    port map (
      a => LPM_q_ivl_21826,
      b => LPM_q_ivl_21835,
      c => LPM_d0_ivl_21843
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4006
  U3886: xnor_HPC2
    port map (
      a => LPM_q_ivl_21847,
      b => LPM_q_ivl_21854,
      c => LPM_d0_ivl_21862
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4007
  U3887: xnor_HPC2
    port map (
      a => LPM_q_ivl_21866,
      b => LPM_q_ivl_21873,
      c => LPM_d0_ivl_21885
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4008
  U3888: xnor_HPC2
    port map (
      a => LPM_q_ivl_21889,
      b => LPM_q_ivl_21896,
      c => LPM_d0_ivl_21904
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4009
  U3889: xnor_HPC2
    port map (
      a => LPM_q_ivl_21908,
      b => LPM_q_ivl_21915,
      c => LPM_d0_ivl_21927
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4010
  U3890: xnor_HPC2
    port map (
      a => LPM_q_ivl_21931,
      b => LPM_q_ivl_21938,
      c => LPM_d0_ivl_21946
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4011
  U3891: xnor_HPC2
    port map (
      a => LPM_q_ivl_21954,
      b => LPM_q_ivl_21961,
      c => LPM_d0_ivl_21969
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4012
  U3892: xnor_HPC2
    port map (
      a => LPM_q_ivl_21973,
      b => LPM_q_ivl_21980,
      c => LPM_d0_ivl_21992
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4013
  U3893: xnor_HPC2
    port map (
      a => LPM_q_ivl_21996,
      b => LPM_q_ivl_22003,
      c => LPM_d0_ivl_22011
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4014
  U3894: xnor_HPC2
    port map (
      a => LPM_q_ivl_22015,
      b => LPM_q_ivl_22022,
      c => LPM_d0_ivl_22034
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4015
  U3895: xnor_HPC2
    port map (
      a => LPM_q_ivl_22038,
      b => LPM_q_ivl_22045,
      c => LPM_d0_ivl_22053
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4016
  U3896: xnor_HPC2
    port map (
      a => LPM_q_ivl_22057,
      b => LPM_q_ivl_22064,
      c => LPM_d0_ivl_22076
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4017
  U3897: xnor_HPC2
    port map (
      a => LPM_q_ivl_22080,
      b => LPM_q_ivl_22087,
      c => LPM_d0_ivl_22095
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4018
  U3898: xor_HPC2
    port map (
      a => LPM_q_ivl_22101,
      b => LPM_q_ivl_22112,
      c => LPM_d0_ivl_22120
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4019
  U3899: xnor_HPC2
    port map (
      a => LPM_q_ivl_22124,
      b => LPM_q_ivl_22131,
      c => LPM_d0_ivl_22139
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4020
  U3900: xnor_HPC2
    port map (
      a => LPM_q_ivl_22143,
      b => LPM_q_ivl_22150,
      c => LPM_d0_ivl_22162
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4021
  U3901: xnor_HPC2
    port map (
      a => LPM_q_ivl_22166,
      b => LPM_q_ivl_22173,
      c => LPM_d0_ivl_22181
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4022
  U3902: xnor_HPC2
    port map (
      a => LPM_q_ivl_22185,
      b => LPM_q_ivl_22192,
      c => LPM_d0_ivl_22204
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4023
  U3903: xnor_HPC2
    port map (
      a => LPM_q_ivl_22208,
      b => LPM_q_ivl_22215,
      c => LPM_d0_ivl_22223
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4024
  U3904: xnor_HPC2
    port map (
      a => LPM_q_ivl_22227,
      b => LPM_q_ivl_22234,
      c => LPM_d0_ivl_22246
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4025
  U3905: xnor_HPC2
    port map (
      a => LPM_q_ivl_22250,
      b => LPM_q_ivl_22257,
      c => LPM_d0_ivl_22265
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4026
  U3906: xor_HPC2
    port map (
      a => LPM_q_ivl_22271,
      b => LPM_q_ivl_22282,
      c => LPM_d0_ivl_22290
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4027
  U3907: xnor_HPC2
    port map (
      a => LPM_q_ivl_22298,
      b => LPM_q_ivl_22305,
      c => LPM_d0_ivl_22313
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4028
  U3908: xnor_HPC2
    port map (
      a => LPM_q_ivl_22317,
      b => LPM_q_ivl_22324,
      c => LPM_d0_ivl_22332
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4029
  U3909: xnor_HPC2
    port map (
      a => LPM_q_ivl_22336,
      b => LPM_q_ivl_22343,
      c => LPM_d0_ivl_22355
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4030
  U3910: xnor_HPC2
    port map (
      a => LPM_q_ivl_22359,
      b => LPM_q_ivl_22366,
      c => LPM_d0_ivl_22374
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4031
  U3911: xnor_HPC2
    port map (
      a => LPM_q_ivl_22378,
      b => LPM_q_ivl_22385,
      c => LPM_d0_ivl_22397
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4032
  U3912: xnor_HPC2
    port map (
      a => LPM_q_ivl_22401,
      b => LPM_q_ivl_22408,
      c => LPM_d0_ivl_22416
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4033
  U3913: xnor_HPC2
    port map (
      a => LPM_q_ivl_22420,
      b => LPM_q_ivl_22427,
      c => LPM_d0_ivl_22439
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4034
  U3914: xnor_HPC2
    port map (
      a => LPM_q_ivl_22443,
      b => LPM_q_ivl_22450,
      c => LPM_d0_ivl_22458
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4035
  U3915: xor_HPC2
    port map (
      a => LPM_q_ivl_22464,
      b => LPM_q_ivl_22475,
      c => LPM_d0_ivl_22483
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4036
  U3916: xnor_HPC2
    port map (
      a => LPM_q_ivl_22487,
      b => LPM_q_ivl_22494,
      c => LPM_d0_ivl_22502
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4037
  U3917: xnor_HPC2
    port map (
      a => LPM_q_ivl_22506,
      b => LPM_q_ivl_22513,
      c => LPM_d0_ivl_22525
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4038
  U3918: xnor_HPC2
    port map (
      a => LPM_q_ivl_22529,
      b => LPM_q_ivl_22536,
      c => LPM_d0_ivl_22544
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4039
  U3919: xnor_HPC2
    port map (
      a => LPM_q_ivl_22548,
      b => LPM_q_ivl_22555,
      c => LPM_d0_ivl_22567
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4040
  U3920: xnor_HPC2
    port map (
      a => LPM_q_ivl_22571,
      b => LPM_q_ivl_22578,
      c => LPM_d0_ivl_22586
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4041
  U3921: xor_HPC2
    port map (
      a => LPM_q_ivl_22592,
      b => LPM_q_ivl_22603,
      c => LPM_d0_ivl_22611
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4042
  U3922: xnor_HPC2
    port map (
      a => LPM_q_ivl_22619,
      b => LPM_q_ivl_22626,
      c => LPM_d0_ivl_22634
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4043
  U3923: xnor_HPC2
    port map (
      a => LPM_q_ivl_22638,
      b => LPM_q_ivl_22645,
      c => LPM_d0_ivl_22653
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4044
  U3924: xnor_HPC2
    port map (
      a => LPM_q_ivl_22657,
      b => LPM_q_ivl_22664,
      c => LPM_d0_ivl_22676
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4045
  U3925: xnor_HPC2
    port map (
      a => LPM_q_ivl_22680,
      b => LPM_q_ivl_22687,
      c => LPM_d0_ivl_22695
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4046
  U3926: xnor_HPC2
    port map (
      a => LPM_q_ivl_22699,
      b => LPM_q_ivl_22706,
      c => LPM_d0_ivl_22718
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4047
  U3927: xnor_HPC2
    port map (
      a => LPM_q_ivl_22722,
      b => LPM_q_ivl_22729,
      c => LPM_d0_ivl_22737
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4048
  U3928: xnor_HPC2
    port map (
      a => LPM_q_ivl_22741,
      b => LPM_q_ivl_22748,
      c => LPM_d0_ivl_22756
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4049
  U3929: xnor_HPC2
    port map (
      a => LPM_q_ivl_22764,
      b => LPM_q_ivl_22773,
      c => LPM_d0_ivl_22781
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4050
  U3930: xnor_HPC2
    port map (
      a => LPM_q_ivl_22785,
      b => LPM_q_ivl_22792,
      c => LPM_d0_ivl_22800
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4051
  U3931: xnor_HPC2
    port map (
      a => LPM_q_ivl_22804,
      b => LPM_q_ivl_22811,
      c => LPM_d0_ivl_22823
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4052
  U3932: xnor_HPC2
    port map (
      a => LPM_q_ivl_22827,
      b => LPM_q_ivl_22834,
      c => LPM_d0_ivl_22842
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4053
  U3933: xnor_HPC2
    port map (
      a => LPM_q_ivl_22846,
      b => LPM_q_ivl_22853,
      c => LPM_d0_ivl_22865
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4054
  U3934: xnor_HPC2
    port map (
      a => LPM_q_ivl_22869,
      b => LPM_q_ivl_22876,
      c => LPM_d0_ivl_22884
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4055
  U3935: xnor_HPC2
    port map (
      a => LPM_q_ivl_22892,
      b => LPM_q_ivl_22899,
      c => LPM_d0_ivl_22907
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4056
  U3936: xnor_HPC2
    port map (
      a => LPM_q_ivl_22911,
      b => LPM_q_ivl_22918,
      c => LPM_d0_ivl_22930
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4057
  U3937: xnor_HPC2
    port map (
      a => LPM_q_ivl_22934,
      b => LPM_q_ivl_22941,
      c => LPM_d0_ivl_22949
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4058
  U3938: xnor_HPC2
    port map (
      a => LPM_q_ivl_22953,
      b => LPM_q_ivl_22960,
      c => LPM_d0_ivl_22972
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4059
  U3939: xnor_HPC2
    port map (
      a => LPM_q_ivl_22976,
      b => LPM_q_ivl_22983,
      c => LPM_d0_ivl_22991
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4060
  U3940: xor_HPC2
    port map (
      a => LPM_q_ivl_22997,
      b => LPM_q_ivl_23008,
      c => LPM_d0_ivl_23016
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4061
  U3941: xnor_HPC2
    port map (
      a => LPM_q_ivl_23020,
      b => LPM_q_ivl_23027,
      c => LPM_d0_ivl_23035
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4062
  U3942: xnor_HPC2
    port map (
      a => LPM_q_ivl_23039,
      b => LPM_q_ivl_23046,
      c => LPM_d0_ivl_23058
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4063
  U3943: xnor_HPC2
    port map (
      a => LPM_q_ivl_23062,
      b => LPM_q_ivl_23069,
      c => LPM_d0_ivl_23077
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4064
  U3944: xnor_HPC2
    port map (
      a => LPM_q_ivl_23081,
      b => LPM_q_ivl_23088,
      c => LPM_d0_ivl_23100
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4065
  U3945: xnor_HPC2
    port map (
      a => LPM_q_ivl_23104,
      b => LPM_q_ivl_23111,
      c => LPM_d0_ivl_23119
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4066
  U3946: xnor_HPC2
    port map (
      a => LPM_q_ivl_23123,
      b => LPM_q_ivl_23130,
      c => LPM_d0_ivl_23142
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4067
  U3947: xnor_HPC2
    port map (
      a => LPM_q_ivl_23146,
      b => LPM_q_ivl_23153,
      c => LPM_d0_ivl_23161
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4068
  U3948: xor_HPC2
    port map (
      a => LPM_q_ivl_23167,
      b => LPM_q_ivl_23174,
      c => LPM_d0_ivl_23182
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3084
  U3949: xnor_HPC2
    port map (
      a => LPM_q_ivl_4151,
      b => LPM_q_ivl_4162,
      c => LPM_d0_ivl_4170
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4069
  U3950: xnor_HPC2
    port map (
      a => LPM_q_ivl_23186,
      b => LPM_q_ivl_23193,
      c => LPM_d0_ivl_23201
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4070
  U3951: xnor_HPC2
    port map (
      a => LPM_q_ivl_23205,
      b => LPM_q_ivl_23212,
      c => LPM_d0_ivl_23224
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4071
  U3952: xnor_HPC2
    port map (
      a => LPM_q_ivl_23228,
      b => LPM_q_ivl_23235,
      c => LPM_d0_ivl_23243
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4072
  U3953: xnor_HPC2
    port map (
      a => LPM_q_ivl_23247,
      b => LPM_q_ivl_23254,
      c => LPM_d0_ivl_23266
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4073
  U3954: xnor_HPC2
    port map (
      a => LPM_q_ivl_23270,
      b => LPM_q_ivl_23277,
      c => LPM_d0_ivl_23285
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4074
  U3955: xor_HPC2
    port map (
      a => LPM_q_ivl_23291,
      b => LPM_q_ivl_23302,
      c => LPM_d0_ivl_23310
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4075
  U3956: xnor_HPC2
    port map (
      a => LPM_q_ivl_23314,
      b => LPM_q_ivl_23321,
      c => LPM_d0_ivl_23329
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4076
  U3957: xnor_HPC2
    port map (
      a => LPM_q_ivl_23333,
      b => LPM_q_ivl_23340,
      c => LPM_d0_ivl_23352
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4077
  U3958: xnor_HPC2
    port map (
      a => LPM_q_ivl_23356,
      b => LPM_q_ivl_23363,
      c => LPM_d0_ivl_23371
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4078
  U3959: xnor_HPC2
    port map (
      a => LPM_q_ivl_23375,
      b => LPM_q_ivl_23382,
      c => LPM_d0_ivl_23394
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4079
  U3960: xnor_HPC2
    port map (
      a => LPM_q_ivl_23398,
      b => LPM_q_ivl_23405,
      c => LPM_d0_ivl_23413
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4080
  U3961: xnor_HPC2
    port map (
      a => LPM_q_ivl_23417,
      b => LPM_q_ivl_23424,
      c => LPM_d0_ivl_23436
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4081
  U3962: xnor_HPC2
    port map (
      a => LPM_q_ivl_23440,
      b => LPM_q_ivl_23447,
      c => LPM_d0_ivl_23455
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4082
  U3963: xor_HPC2
    port map (
      a => LPM_q_ivl_23461,
      b => LPM_q_ivl_23472,
      c => LPM_d0_ivl_23480
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4083
  U3964: xnor_HPC2
    port map (
      a => LPM_q_ivl_23488,
      b => LPM_q_ivl_23495,
      c => LPM_d0_ivl_23503
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4084
  U3965: xnor_HPC2
    port map (
      a => LPM_q_ivl_23507,
      b => LPM_q_ivl_23514,
      c => LPM_d0_ivl_23522
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4085
  U3966: xnor_HPC2
    port map (
      a => LPM_q_ivl_23526,
      b => LPM_q_ivl_23533,
      c => LPM_d0_ivl_23545
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4086
  U3967: xnor_HPC2
    port map (
      a => LPM_q_ivl_23549,
      b => LPM_q_ivl_23556,
      c => LPM_d0_ivl_23564
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4087
  U3968: xnor_HPC2
    port map (
      a => LPM_q_ivl_23568,
      b => LPM_q_ivl_23575,
      c => LPM_d0_ivl_23587
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4088
  U3969: xnor_HPC2
    port map (
      a => LPM_q_ivl_23591,
      b => LPM_q_ivl_23598,
      c => LPM_d0_ivl_23606
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4089
  U3970: xnor_HPC2
    port map (
      a => LPM_q_ivl_23610,
      b => LPM_q_ivl_23617,
      c => LPM_d0_ivl_23629
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4090
  U3971: xnor_HPC2
    port map (
      a => LPM_q_ivl_23633,
      b => LPM_q_ivl_23640,
      c => LPM_d0_ivl_23648
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4091
  U3972: xnor_HPC2
    port map (
      a => LPM_q_ivl_23656,
      b => LPM_q_ivl_23665,
      c => LPM_d0_ivl_23673
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4092
  U3973: xnor_HPC2
    port map (
      a => LPM_q_ivl_23677,
      b => LPM_q_ivl_23684,
      c => LPM_d0_ivl_23692
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4093
  U3974: xnor_HPC2
    port map (
      a => LPM_q_ivl_23696,
      b => LPM_q_ivl_23703,
      c => LPM_d0_ivl_23715
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4094
  U3975: xnor_HPC2
    port map (
      a => LPM_q_ivl_23719,
      b => LPM_q_ivl_23726,
      c => LPM_d0_ivl_23734
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4095
  U3976: xnor_HPC2
    port map (
      a => LPM_q_ivl_23738,
      b => LPM_q_ivl_23745,
      c => LPM_d0_ivl_23757
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4096
  U3977: xnor_HPC2
    port map (
      a => LPM_q_ivl_23761,
      b => LPM_q_ivl_23768,
      c => LPM_d0_ivl_23776
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4097
  U3978: xnor_HPC2
    port map (
      a => LPM_q_ivl_23780,
      b => LPM_q_ivl_23787,
      c => LPM_d0_ivl_23799
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4098
  U3979: xnor_HPC2
    port map (
      a => LPM_q_ivl_23803,
      b => LPM_q_ivl_23810,
      c => LPM_d0_ivl_23818
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4099
  U3980: xnor_HPC2
    port map (
      a => LPM_q_ivl_23826,
      b => LPM_q_ivl_23833,
      c => LPM_d0_ivl_23841
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4100
  U3981: xnor_HPC2
    port map (
      a => LPM_q_ivl_23845,
      b => LPM_q_ivl_23852,
      c => LPM_d0_ivl_23864
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4101
  U3982: xnor_HPC2
    port map (
      a => LPM_q_ivl_23868,
      b => LPM_q_ivl_23875,
      c => LPM_d0_ivl_23883
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4102
  U3983: xnor_HPC2
    port map (
      a => LPM_q_ivl_23887,
      b => LPM_q_ivl_23894,
      c => LPM_d0_ivl_23906
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4103
  U3984: xnor_HPC2
    port map (
      a => LPM_q_ivl_23910,
      b => LPM_q_ivl_23917,
      c => LPM_d0_ivl_23925
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4104
  U3985: xnor_HPC2
    port map (
      a => LPM_q_ivl_23929,
      b => LPM_q_ivl_23936,
      c => LPM_d0_ivl_23948
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4105
  U3986: xnor_HPC2
    port map (
      a => LPM_q_ivl_23952,
      b => LPM_q_ivl_23959,
      c => LPM_d0_ivl_23967
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4106
  U3987: xor_HPC2
    port map (
      a => LPM_q_ivl_23973,
      b => LPM_q_ivl_23984,
      c => LPM_d0_ivl_23992
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4107
  U3988: xnor_HPC2
    port map (
      a => LPM_q_ivl_23996,
      b => LPM_q_ivl_24003,
      c => LPM_d0_ivl_24011
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4108
  U3989: xnor_HPC2
    port map (
      a => LPM_q_ivl_24015,
      b => LPM_q_ivl_24022,
      c => LPM_d0_ivl_24034
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4109
  U3990: xnor_HPC2
    port map (
      a => LPM_q_ivl_24038,
      b => LPM_q_ivl_24045,
      c => LPM_d0_ivl_24053
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4110
  U3991: xnor_HPC2
    port map (
      a => LPM_q_ivl_24057,
      b => LPM_q_ivl_24064,
      c => LPM_d0_ivl_24076
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4111
  U3992: xnor_HPC2
    port map (
      a => LPM_q_ivl_24080,
      b => LPM_q_ivl_24087,
      c => LPM_d0_ivl_24095
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4112
  U3993: xor_HPC2
    port map (
      a => LPM_q_ivl_24101,
      b => LPM_q_ivl_24112,
      c => LPM_d0_ivl_24120
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4113
  U3994: xnor_HPC2
    port map (
      a => LPM_q_ivl_24128,
      b => LPM_q_ivl_24135,
      c => LPM_d0_ivl_24143
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4114
  U3995: xnor_HPC2
    port map (
      a => LPM_q_ivl_24147,
      b => LPM_q_ivl_24154,
      c => LPM_d0_ivl_24162
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4115
  U3996: xnor_HPC2
    port map (
      a => LPM_q_ivl_24166,
      b => LPM_q_ivl_24173,
      c => LPM_d0_ivl_24185
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4116
  U3997: xnor_HPC2
    port map (
      a => LPM_q_ivl_24189,
      b => LPM_q_ivl_24196,
      c => LPM_d0_ivl_24204
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4117
  U3998: xnor_HPC2
    port map (
      a => LPM_q_ivl_24208,
      b => LPM_q_ivl_24215,
      c => LPM_d0_ivl_24227
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4118
  U3999: xnor_HPC2
    port map (
      a => LPM_q_ivl_24231,
      b => LPM_q_ivl_24238,
      c => LPM_d0_ivl_24246
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4119
  U4000: xnor_HPC2
    port map (
      a => LPM_q_ivl_24254,
      b => LPM_q_ivl_24263,
      c => LPM_d0_ivl_24271
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4120
  U4001: xnor_HPC2
    port map (
      a => LPM_q_ivl_24275,
      b => LPM_q_ivl_24282,
      c => LPM_d0_ivl_24290
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4121
  U4002: xnor_HPC2
    port map (
      a => LPM_q_ivl_24294,
      b => LPM_q_ivl_24301,
      c => LPM_d0_ivl_24313
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4122
  U4003: xnor_HPC2
    port map (
      a => LPM_q_ivl_24317,
      b => LPM_q_ivl_24324,
      c => LPM_d0_ivl_24332
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4123
  U4004: xnor_HPC2
    port map (
      a => LPM_q_ivl_24336,
      b => LPM_q_ivl_24343,
      c => LPM_d0_ivl_24355
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4124
  U4005: xnor_HPC2
    port map (
      a => LPM_q_ivl_24359,
      b => LPM_q_ivl_24366,
      c => LPM_d0_ivl_24374
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4125
  U4006: xnor_HPC2
    port map (
      a => LPM_q_ivl_24378,
      b => LPM_q_ivl_24385,
      c => LPM_d0_ivl_24397
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4126
  U4007: xnor_HPC2
    port map (
      a => LPM_q_ivl_24401,
      b => LPM_q_ivl_24408,
      c => LPM_d0_ivl_24416
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4127
  U4008: xnor_HPC2
    port map (
      a => LPM_q_ivl_24424,
      b => LPM_q_ivl_24431,
      c => LPM_d0_ivl_24439
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4128
  U4009: xnor_HPC2
    port map (
      a => LPM_q_ivl_24443,
      b => LPM_q_ivl_24450,
      c => LPM_d0_ivl_24462
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4129
  U4010: xnor_HPC2
    port map (
      a => LPM_q_ivl_24466,
      b => LPM_q_ivl_24473,
      c => LPM_d0_ivl_24481
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4130
  U4011: xnor_HPC2
    port map (
      a => LPM_q_ivl_24485,
      b => LPM_q_ivl_24492,
      c => LPM_d0_ivl_24504
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4131
  U4012: xnor_HPC2
    port map (
      a => LPM_q_ivl_24508,
      b => LPM_q_ivl_24515,
      c => LPM_d0_ivl_24523
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4132
  U4013: xor_HPC2
    port map (
      a => LPM_q_ivl_24529,
      b => LPM_q_ivl_24540,
      c => LPM_d0_ivl_24548
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4133
  U4014: xnor_HPC2
    port map (
      a => LPM_q_ivl_24552,
      b => LPM_q_ivl_24559,
      c => LPM_d0_ivl_24567
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4134
  U4015: xnor_HPC2
    port map (
      a => LPM_q_ivl_24571,
      b => LPM_q_ivl_24578,
      c => LPM_d0_ivl_24590
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4135
  U4016: xnor_HPC2
    port map (
      a => LPM_q_ivl_24594,
      b => LPM_q_ivl_24601,
      c => LPM_d0_ivl_24609
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4136
  U4017: xnor_HPC2
    port map (
      a => LPM_q_ivl_24613,
      b => LPM_q_ivl_24620,
      c => LPM_d0_ivl_24632
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4137
  U4018: xnor_HPC2
    port map (
      a => LPM_q_ivl_24636,
      b => LPM_q_ivl_24643,
      c => LPM_d0_ivl_24651
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4138
  U4019: xor_HPC2
    port map (
      a => LPM_q_ivl_24657,
      b => LPM_q_ivl_24668,
      c => LPM_d0_ivl_24676
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4139
  U4020: xnor_HPC2
    port map (
      a => LPM_q_ivl_24684,
      b => LPM_q_ivl_24691,
      c => LPM_d0_ivl_24699
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4140
  U4021: xnor_HPC2
    port map (
      a => LPM_q_ivl_24703,
      b => LPM_q_ivl_24710,
      c => LPM_d0_ivl_24718
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4141
  U4022: xnor_HPC2
    port map (
      a => LPM_q_ivl_24722,
      b => LPM_q_ivl_24729,
      c => LPM_d0_ivl_24741
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4142
  U4023: xnor_HPC2
    port map (
      a => LPM_q_ivl_24745,
      b => LPM_q_ivl_24752,
      c => LPM_d0_ivl_24760
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4143
  U4024: xnor_HPC2
    port map (
      a => LPM_q_ivl_24764,
      b => LPM_q_ivl_24771,
      c => LPM_d0_ivl_24783
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4144
  U4025: xnor_HPC2
    port map (
      a => LPM_q_ivl_24787,
      b => LPM_q_ivl_24794,
      c => LPM_d0_ivl_24802
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4145
  U4026: xor_HPC2
    port map (
      a => LPM_q_ivl_24808,
      b => LPM_q_ivl_24819,
      c => LPM_d0_ivl_24827
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4146
  U4027: xnor_HPC2
    port map (
      a => LPM_q_ivl_24831,
      b => LPM_q_ivl_24838,
      c => LPM_d0_ivl_24846
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4147
  U4028: xnor_HPC2
    port map (
      a => LPM_q_ivl_24850,
      b => LPM_q_ivl_24857,
      c => LPM_d0_ivl_24869
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4148
  U4029: xnor_HPC2
    port map (
      a => LPM_q_ivl_24873,
      b => LPM_q_ivl_24880,
      c => LPM_d0_ivl_24888
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4149
  U4030: xnor_HPC2
    port map (
      a => LPM_q_ivl_24892,
      b => LPM_q_ivl_24899,
      c => LPM_d0_ivl_24911
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4150
  U4031: xnor_HPC2
    port map (
      a => LPM_q_ivl_24915,
      b => LPM_q_ivl_24922,
      c => LPM_d0_ivl_24930
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4151
  U4032: xnor_HPC2
    port map (
      a => LPM_q_ivl_24934,
      b => LPM_q_ivl_24941,
      c => LPM_d0_ivl_24953
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4152
  U4033: xnor_HPC2
    port map (
      a => LPM_q_ivl_24957,
      b => LPM_q_ivl_24964,
      c => LPM_d0_ivl_24972
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4153
  U4034: xor_HPC2
    port map (
      a => LPM_q_ivl_24978,
      b => LPM_q_ivl_24989,
      c => LPM_d0_ivl_24997
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4154
  U4035: xnor_HPC2
    port map (
      a => LPM_q_ivl_25005,
      b => LPM_q_ivl_25012,
      c => LPM_d0_ivl_25020
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4155
  U4036: xnor_HPC2
    port map (
      a => LPM_q_ivl_25024,
      b => LPM_q_ivl_25031,
      c => LPM_d0_ivl_25039
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4156
  U4037: xnor_HPC2
    port map (
      a => LPM_q_ivl_25043,
      b => LPM_q_ivl_25050,
      c => LPM_d0_ivl_25062
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4157
  U4038: xnor_HPC2
    port map (
      a => LPM_q_ivl_25066,
      b => LPM_q_ivl_25073,
      c => LPM_d0_ivl_25081
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4158
  U4039: xnor_HPC2
    port map (
      a => LPM_q_ivl_25085,
      b => LPM_q_ivl_25092,
      c => LPM_d0_ivl_25104
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4159
  U4040: xnor_HPC2
    port map (
      a => LPM_q_ivl_25108,
      b => LPM_q_ivl_25115,
      c => LPM_d0_ivl_25123
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4160
  U4041: xnor_HPC2
    port map (
      a => LPM_q_ivl_25127,
      b => LPM_q_ivl_25134,
      c => LPM_d0_ivl_25146
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4161
  U4042: xnor_HPC2
    port map (
      a => LPM_q_ivl_25150,
      b => LPM_q_ivl_25157,
      c => LPM_d0_ivl_25165
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4162
  U4043: xnor_HPC2
    port map (
      a => LPM_q_ivl_25173,
      b => LPM_q_ivl_25182,
      c => LPM_d0_ivl_25190
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4163
  U4044: xnor_HPC2
    port map (
      a => LPM_q_ivl_25194,
      b => LPM_q_ivl_25201,
      c => LPM_d0_ivl_25209
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4164
  U4045: xnor_HPC2
    port map (
      a => LPM_q_ivl_25213,
      b => LPM_q_ivl_25220,
      c => LPM_d0_ivl_25232
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4165
  U4046: xnor_HPC2
    port map (
      a => LPM_q_ivl_25236,
      b => LPM_q_ivl_25243,
      c => LPM_d0_ivl_25251
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4166
  U4047: xnor_HPC2
    port map (
      a => LPM_q_ivl_25255,
      b => LPM_q_ivl_25262,
      c => LPM_d0_ivl_25274
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4167
  U4048: xnor_HPC2
    port map (
      a => LPM_q_ivl_25278,
      b => LPM_q_ivl_25285,
      c => LPM_d0_ivl_25293
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4168
  U4049: xnor_HPC2
    port map (
      a => LPM_q_ivl_25297,
      b => LPM_q_ivl_25304,
      c => LPM_d0_ivl_25316
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4169
  U4050: xnor_HPC2
    port map (
      a => LPM_q_ivl_25320,
      b => LPM_q_ivl_25327,
      c => LPM_d0_ivl_25335
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4170
  U4051: xnor_HPC2
    port map (
      a => LPM_q_ivl_25343,
      b => LPM_q_ivl_25350,
      c => LPM_d0_ivl_25358
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4171
  U4052: xnor_HPC2
    port map (
      a => LPM_q_ivl_25362,
      b => LPM_q_ivl_25369,
      c => LPM_d0_ivl_25381
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4172
  U4053: xnor_HPC2
    port map (
      a => LPM_q_ivl_25385,
      b => LPM_q_ivl_25392,
      c => LPM_d0_ivl_25400
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4173
  U4054: xnor_HPC2
    port map (
      a => LPM_q_ivl_25404,
      b => LPM_q_ivl_25411,
      c => LPM_d0_ivl_25423
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4174
  U4055: xnor_HPC2
    port map (
      a => LPM_q_ivl_25427,
      b => LPM_q_ivl_25434,
      c => LPM_d0_ivl_25442
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4175
  U4056: xnor_HPC2
    port map (
      a => LPM_q_ivl_25446,
      b => LPM_q_ivl_25453,
      c => LPM_d0_ivl_25465
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3085
  U4057: xor_HPC2
    port map (
      a => LPM_q_ivl_4178,
      b => LPM_q_ivl_4189,
      c => LPM_d0_ivl_4197
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3086
  U4058: xor_HPC2
    port map (
      a => LPM_q_ivl_4205,
      b => LPM_q_ivl_4216,
      c => LPM_d0_ivl_4224
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3087
  U4059: xor_HPC2
    port map (
      a => LPM_q_ivl_4232,
      b => LPM_q_ivl_4243,
      c => LPM_d0_ivl_4251
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4176
  U4060: xor_HPC2
    port map (
      a => LPM_q_ivl_25469,
      b => LPM_q_ivl_25478,
      c => LPM_d0_ivl_25486
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4177
  U4061: xnor_HPC2
    port map (
      a => LPM_q_ivl_25492,
      b => LPM_q_ivl_25503,
      c => LPM_d0_ivl_25511
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4178
  U4062: xnor_HPC2
    port map (
      a => LPM_q_ivl_25515,
      b => LPM_q_ivl_25522,
      c => LPM_d0_ivl_25530
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4179
  U4063: xor_HPC2
    port map (
      a => LPM_q_ivl_25534,
      b => LPM_q_ivl_25543,
      c => LPM_d0_ivl_25551
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4180
  U4064: xor_HPC2
    port map (
      a => LPM_q_ivl_25557,
      b => LPM_q_ivl_25568,
      c => LPM_d0_ivl_25576
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4181
  U4065: xnor_HPC2
    port map (
      a => LPM_q_ivl_25580,
      b => LPM_q_ivl_25587,
      c => LPM_d0_ivl_25595
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4182
  U4066: xnor_HPC2
    port map (
      a => LPM_q_ivl_25599,
      b => LPM_q_ivl_25606,
      c => LPM_d0_ivl_25614
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4183
  U4067: xor_HPC2
    port map (
      a => LPM_q_ivl_25618,
      b => LPM_q_ivl_25627,
      c => LPM_d0_ivl_25635
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4184
  U4068: xor_HPC2
    port map (
      a => LPM_q_ivl_25641,
      b => LPM_q_ivl_25652,
      c => LPM_d0_ivl_25660
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4185
  U4069: xnor_HPC2
    port map (
      a => LPM_q_ivl_25664,
      b => LPM_q_ivl_25671,
      c => LPM_d0_ivl_25679
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4186
  U4070: xnor_HPC2
    port map (
      a => LPM_q_ivl_25683,
      b => LPM_q_ivl_25690,
      c => LPM_d0_ivl_25702
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3088
  U4071: xor_HPC2
    port map (
      a => LPM_q_ivl_4259,
      b => LPM_q_ivl_4270,
      c => LPM_d0_ivl_4278
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3089
  U4072: xor_HPC2
    port map (
      a => LPM_q_ivl_4286,
      b => LPM_q_ivl_4297,
      c => LPM_d0_ivl_4305
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3090
  U4073: xor_HPC2
    port map (
      a => LPM_q_ivl_4313,
      b => LPM_q_ivl_4324,
      c => LPM_d0_ivl_4332
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4187
  U4074: xor_HPC2
    port map (
      a => LPM_q_ivl_25706,
      b => LPM_q_ivl_25715,
      c => LPM_d0_ivl_25723
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4188
  U4075: xnor_HPC2
    port map (
      a => LPM_q_ivl_25729,
      b => LPM_q_ivl_25740,
      c => LPM_d0_ivl_25748
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4189
  U4076: xnor_HPC2
    port map (
      a => LPM_q_ivl_25752,
      b => LPM_q_ivl_25759,
      c => LPM_d0_ivl_25767
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4190
  U4077: xor_HPC2
    port map (
      a => LPM_q_ivl_25771,
      b => LPM_q_ivl_25780,
      c => LPM_d0_ivl_25788
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4191
  U4078: xor_HPC2
    port map (
      a => LPM_q_ivl_25794,
      b => LPM_q_ivl_25805,
      c => LPM_d0_ivl_25813
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4192
  U4079: xnor_HPC2
    port map (
      a => LPM_q_ivl_25817,
      b => LPM_q_ivl_25824,
      c => LPM_d0_ivl_25832
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4193
  U4080: xnor_HPC2
    port map (
      a => LPM_q_ivl_25836,
      b => LPM_q_ivl_25843,
      c => LPM_d0_ivl_25851
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4194
  U4081: xor_HPC2
    port map (
      a => LPM_q_ivl_25855,
      b => LPM_q_ivl_25864,
      c => LPM_d0_ivl_25872
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4195
  U4082: xor_HPC2
    port map (
      a => LPM_q_ivl_25878,
      b => LPM_q_ivl_25889,
      c => LPM_d0_ivl_25897
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4196
  U4083: xnor_HPC2
    port map (
      a => LPM_q_ivl_25901,
      b => LPM_q_ivl_25908,
      c => LPM_d0_ivl_25916
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4197
  U4084: xnor_HPC2
    port map (
      a => LPM_q_ivl_25920,
      b => LPM_q_ivl_25927,
      c => LPM_d0_ivl_25939
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3091
  U4085: xor_HPC2
    port map (
      a => LPM_q_ivl_4340,
      b => LPM_q_ivl_4351,
      c => LPM_d0_ivl_4359
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3092
  U4086: xor_HPC2
    port map (
      a => LPM_q_ivl_4367,
      b => LPM_q_ivl_4378,
      c => LPM_d0_ivl_4386
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3093
  U4087: xor_HPC2
    port map (
      a => LPM_q_ivl_4394,
      b => LPM_q_ivl_4405,
      c => LPM_d0_ivl_4413
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4198
  U4088: xor_HPC2
    port map (
      a => LPM_q_ivl_25943,
      b => LPM_q_ivl_25952,
      c => LPM_d0_ivl_25960
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4199
  U4089: xnor_HPC2
    port map (
      a => LPM_q_ivl_25966,
      b => LPM_q_ivl_25977,
      c => LPM_d0_ivl_25985
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4200
  U4090: xnor_HPC2
    port map (
      a => LPM_q_ivl_25989,
      b => LPM_q_ivl_25996,
      c => LPM_d0_ivl_26004
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4201
  U4091: xor_HPC2
    port map (
      a => LPM_q_ivl_26008,
      b => LPM_q_ivl_26017,
      c => LPM_d0_ivl_26025
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4202
  U4092: xnor_HPC2
    port map (
      a => LPM_q_ivl_26031,
      b => LPM_q_ivl_26042,
      c => LPM_d0_ivl_26050
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4203
  U4093: xnor_HPC2
    port map (
      a => LPM_q_ivl_26054,
      b => LPM_q_ivl_26061,
      c => LPM_d0_ivl_26069
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4204
  U4094: xor_HPC2
    port map (
      a => LPM_q_ivl_26073,
      b => LPM_q_ivl_26082,
      c => LPM_d0_ivl_26090
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4205
  U4095: xnor_HPC2
    port map (
      a => LPM_q_ivl_26096,
      b => LPM_q_ivl_26107,
      c => LPM_d0_ivl_26115
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4206
  U4096: xnor_HPC2
    port map (
      a => LPM_q_ivl_26119,
      b => LPM_q_ivl_26126,
      c => LPM_d0_ivl_26134
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4207
  U4097: xnor_HPC2
    port map (
      a => LPM_q_ivl_26138,
      b => LPM_q_ivl_26145,
      c => LPM_d0_ivl_26153
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4208
  U4098: xnor_HPC2
    port map (
      a => LPM_q_ivl_26157,
      b => LPM_q_ivl_26164,
      c => LPM_d0_ivl_26176
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3094
  U4099: xor_HPC2
    port map (
      a => LPM_q_ivl_4421,
      b => LPM_q_ivl_4432,
      c => LPM_d0_ivl_4440
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3095
  U4100: xor_HPC2
    port map (
      a => LPM_q_ivl_4448,
      b => LPM_q_ivl_4459,
      c => LPM_d0_ivl_4467
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3096
  U4101: xor_HPC2
    port map (
      a => LPM_q_ivl_4475,
      b => LPM_q_ivl_4486,
      c => LPM_d0_ivl_4494
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4209
  U4102: xor_HPC2
    port map (
      a => LPM_q_ivl_26180,
      b => LPM_q_ivl_26189,
      c => LPM_d0_ivl_26197
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4210
  U4103: xnor_HPC2
    port map (
      a => LPM_q_ivl_26203,
      b => LPM_q_ivl_26214,
      c => LPM_d0_ivl_26222
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4211
  U4104: xnor_HPC2
    port map (
      a => LPM_q_ivl_26226,
      b => LPM_q_ivl_26233,
      c => LPM_d0_ivl_26241
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4212
  U4105: xor_HPC2
    port map (
      a => LPM_q_ivl_26245,
      b => LPM_q_ivl_26254,
      c => LPM_d0_ivl_26262
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4213
  U4106: xnor_HPC2
    port map (
      a => LPM_q_ivl_26268,
      b => LPM_q_ivl_26279,
      c => LPM_d0_ivl_26287
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4214
  U4107: xnor_HPC2
    port map (
      a => LPM_q_ivl_26291,
      b => LPM_q_ivl_26298,
      c => LPM_d0_ivl_26306
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4215
  U4108: xor_HPC2
    port map (
      a => LPM_q_ivl_26310,
      b => LPM_q_ivl_26319,
      c => LPM_d0_ivl_26327
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4216
  U4109: xnor_HPC2
    port map (
      a => LPM_q_ivl_26333,
      b => LPM_q_ivl_26344,
      c => LPM_d0_ivl_26352
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4217
  U4110: xnor_HPC2
    port map (
      a => LPM_q_ivl_26356,
      b => LPM_q_ivl_26363,
      c => LPM_d0_ivl_26371
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4218
  U4111: xnor_HPC2
    port map (
      a => LPM_q_ivl_26375,
      b => LPM_q_ivl_26382,
      c => LPM_d0_ivl_26390
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4219
  U4112: xnor_HPC2
    port map (
      a => LPM_q_ivl_26394,
      b => LPM_q_ivl_26401,
      c => LPM_d0_ivl_26413
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3097
  U4113: xor_HPC2
    port map (
      a => LPM_q_ivl_4502,
      b => LPM_q_ivl_4513,
      c => LPM_d0_ivl_4521
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3098
  U4114: xor_HPC2
    port map (
      a => LPM_q_ivl_4529,
      b => LPM_q_ivl_4540,
      c => LPM_d0_ivl_4548
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3099
  U4115: xor_HPC2
    port map (
      a => LPM_q_ivl_4556,
      b => LPM_q_ivl_4567,
      c => LPM_d0_ivl_4575
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4220
  U4116: xor_HPC2
    port map (
      a => LPM_q_ivl_26417,
      b => LPM_q_ivl_26426,
      c => LPM_d0_ivl_26434
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4221
  U4117: xnor_HPC2
    port map (
      a => LPM_q_ivl_26440,
      b => LPM_q_ivl_26451,
      c => LPM_d0_ivl_26459
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4222
  U4118: xnor_HPC2
    port map (
      a => LPM_q_ivl_26463,
      b => LPM_q_ivl_26470,
      c => LPM_d0_ivl_26478
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4223
  U4119: xor_HPC2
    port map (
      a => LPM_q_ivl_26482,
      b => LPM_q_ivl_26491,
      c => LPM_d0_ivl_26499
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4224
  U4120: xor_HPC2
    port map (
      a => LPM_q_ivl_26505,
      b => LPM_q_ivl_26516,
      c => LPM_d0_ivl_26524
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4225
  U4121: xnor_HPC2
    port map (
      a => LPM_q_ivl_26528,
      b => LPM_q_ivl_26535,
      c => LPM_d0_ivl_26543
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4226
  U4122: xnor_HPC2
    port map (
      a => LPM_q_ivl_26547,
      b => LPM_q_ivl_26554,
      c => LPM_d0_ivl_26562
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4227
  U4123: xor_HPC2
    port map (
      a => LPM_q_ivl_26566,
      b => LPM_q_ivl_26575,
      c => LPM_d0_ivl_26583
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4228
  U4124: xor_HPC2
    port map (
      a => LPM_q_ivl_26589,
      b => LPM_q_ivl_26600,
      c => LPM_d0_ivl_26608
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4229
  U4125: xnor_HPC2
    port map (
      a => LPM_q_ivl_26612,
      b => LPM_q_ivl_26619,
      c => LPM_d0_ivl_26627
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4230
  U4126: xnor_HPC2
    port map (
      a => LPM_q_ivl_26631,
      b => LPM_q_ivl_26638,
      c => LPM_d0_ivl_26650
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3100
  U4127: xor_HPC2
    port map (
      a => LPM_q_ivl_4583,
      b => LPM_q_ivl_4594,
      c => LPM_d0_ivl_4602
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3101
  U4128: xor_HPC2
    port map (
      a => LPM_q_ivl_4610,
      b => LPM_q_ivl_4621,
      c => LPM_d0_ivl_4629
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3102
  U4129: xor_HPC2
    port map (
      a => LPM_q_ivl_4637,
      b => LPM_q_ivl_4648,
      c => LPM_d0_ivl_4656
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4231
  U4130: xor_HPC2
    port map (
      a => LPM_q_ivl_26654,
      b => LPM_q_ivl_26663,
      c => LPM_d0_ivl_26671
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4232
  U4131: xnor_HPC2
    port map (
      a => LPM_q_ivl_26677,
      b => LPM_q_ivl_26688,
      c => LPM_d0_ivl_26696
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4233
  U4132: xnor_HPC2
    port map (
      a => LPM_q_ivl_26700,
      b => LPM_q_ivl_26707,
      c => LPM_d0_ivl_26715
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4234
  U4133: xor_HPC2
    port map (
      a => LPM_q_ivl_26719,
      b => LPM_q_ivl_26728,
      c => LPM_d0_ivl_26736
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4235
  U4134: xnor_HPC2
    port map (
      a => LPM_q_ivl_26742,
      b => LPM_q_ivl_26753,
      c => LPM_d0_ivl_26761
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4236
  U4135: xnor_HPC2
    port map (
      a => LPM_q_ivl_26765,
      b => LPM_q_ivl_26772,
      c => LPM_d0_ivl_26780
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4237
  U4136: xnor_HPC2
    port map (
      a => LPM_q_ivl_26784,
      b => LPM_q_ivl_26791,
      c => LPM_d0_ivl_26799
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4238
  U4137: xor_HPC2
    port map (
      a => LPM_q_ivl_26803,
      b => LPM_q_ivl_26812,
      c => LPM_d0_ivl_26820
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4239
  U4138: xnor_HPC2
    port map (
      a => LPM_q_ivl_26826,
      b => LPM_q_ivl_26837,
      c => LPM_d0_ivl_26845
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4240
  U4139: xnor_HPC2
    port map (
      a => LPM_q_ivl_26849,
      b => LPM_q_ivl_26856,
      c => LPM_d0_ivl_26864
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4241
  U4140: xnor_HPC2
    port map (
      a => LPM_q_ivl_26868,
      b => LPM_q_ivl_26875,
      c => LPM_d0_ivl_26887
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3103
  U4141: xor_HPC2
    port map (
      a => LPM_q_ivl_4664,
      b => LPM_q_ivl_4675,
      c => LPM_d0_ivl_4683
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3104
  U4142: xor_HPC2
    port map (
      a => LPM_q_ivl_4691,
      b => LPM_q_ivl_4702,
      c => LPM_d0_ivl_4710
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3105
  U4143: xor_HPC2
    port map (
      a => LPM_q_ivl_4718,
      b => LPM_q_ivl_4729,
      c => LPM_d0_ivl_4737
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4242
  U4144: xor_HPC2
    port map (
      a => LPM_q_ivl_26891,
      b => LPM_q_ivl_26900,
      c => LPM_d0_ivl_26908
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4243
  U4145: xnor_HPC2
    port map (
      a => LPM_q_ivl_26914,
      b => LPM_q_ivl_26925,
      c => LPM_d0_ivl_26933
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4244
  U4146: xnor_HPC2
    port map (
      a => LPM_q_ivl_26937,
      b => LPM_q_ivl_26944,
      c => LPM_d0_ivl_26952
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4245
  U4147: xor_HPC2
    port map (
      a => LPM_q_ivl_26956,
      b => LPM_q_ivl_26965,
      c => LPM_d0_ivl_26973
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4246
  U4148: xnor_HPC2
    port map (
      a => LPM_q_ivl_26979,
      b => LPM_q_ivl_26990,
      c => LPM_d0_ivl_26998
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4247
  U4149: xnor_HPC2
    port map (
      a => LPM_q_ivl_27002,
      b => LPM_q_ivl_27009,
      c => LPM_d0_ivl_27017
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4248
  U4150: xor_HPC2
    port map (
      a => LPM_q_ivl_27021,
      b => LPM_q_ivl_27030,
      c => LPM_d0_ivl_27038
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4249
  U4151: xnor_HPC2
    port map (
      a => LPM_q_ivl_27044,
      b => LPM_q_ivl_27055,
      c => LPM_d0_ivl_27063
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4250
  U4152: xnor_HPC2
    port map (
      a => LPM_q_ivl_27067,
      b => LPM_q_ivl_27074,
      c => LPM_d0_ivl_27082
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4251
  U4153: xnor_HPC2
    port map (
      a => LPM_q_ivl_27086,
      b => LPM_q_ivl_27093,
      c => LPM_d0_ivl_27101
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4252
  U4154: xnor_HPC2
    port map (
      a => LPM_q_ivl_27105,
      b => LPM_q_ivl_27112,
      c => LPM_d0_ivl_27124
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3106
  U4155: xor_HPC2
    port map (
      a => LPM_q_ivl_4745,
      b => LPM_q_ivl_4756,
      c => LPM_d0_ivl_4764
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3107
  U4156: xor_HPC2
    port map (
      a => LPM_q_ivl_4772,
      b => LPM_q_ivl_4783,
      c => LPM_d0_ivl_4791
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4253
  U4157: xor_HPC2
    port map (
      a => LPM_q_ivl_27128,
      b => LPM_q_ivl_27137,
      c => LPM_d0_ivl_27145
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4254
  U4158: xnor_HPC2
    port map (
      a => LPM_q_ivl_27151,
      b => LPM_q_ivl_27162,
      c => LPM_d0_ivl_27170
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4255
  U4159: xnor_HPC2
    port map (
      a => LPM_q_ivl_27174,
      b => LPM_q_ivl_27181,
      c => LPM_d0_ivl_27189
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4256
  U4160: xnor_HPC2
    port map (
      a => LPM_q_ivl_27193,
      b => LPM_q_ivl_27200,
      c => LPM_d0_ivl_27208
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4257
  U4161: xor_HPC2
    port map (
      a => LPM_q_ivl_27212,
      b => LPM_q_ivl_27221,
      c => LPM_d0_ivl_27229
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4258
  U4162: xor_HPC2
    port map (
      a => LPM_q_ivl_27235,
      b => LPM_q_ivl_27246,
      c => LPM_d0_ivl_27254
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4259
  U4163: xnor_HPC2
    port map (
      a => LPM_q_ivl_27258,
      b => LPM_q_ivl_27265,
      c => LPM_d0_ivl_27273
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4260
  U4164: xnor_HPC2
    port map (
      a => LPM_q_ivl_27277,
      b => LPM_q_ivl_27284,
      c => LPM_d0_ivl_27296
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3108
  U4165: xor_HPC2
    port map (
      a => LPM_q_ivl_4799,
      b => LPM_q_ivl_4810,
      c => LPM_d0_ivl_4818
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3109
  U4166: xor_HPC2
    port map (
      a => LPM_q_ivl_4826,
      b => LPM_q_ivl_4837,
      c => LPM_d0_ivl_4845
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4261
  U4167: xor_HPC2
    port map (
      a => LPM_q_ivl_27300,
      b => LPM_q_ivl_27309,
      c => LPM_d0_ivl_27317
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4262
  U4168: xnor_HPC2
    port map (
      a => LPM_q_ivl_27323,
      b => LPM_q_ivl_27334,
      c => LPM_d0_ivl_27342
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4263
  U4169: xnor_HPC2
    port map (
      a => LPM_q_ivl_27346,
      b => LPM_q_ivl_27353,
      c => LPM_d0_ivl_27361
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4264
  U4170: xnor_HPC2
    port map (
      a => LPM_q_ivl_27365,
      b => LPM_q_ivl_27372,
      c => LPM_d0_ivl_27380
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4265
  U4171: xor_HPC2
    port map (
      a => LPM_q_ivl_27384,
      b => LPM_q_ivl_27393,
      c => LPM_d0_ivl_27401
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4266
  U4172: xor_HPC2
    port map (
      a => LPM_q_ivl_27407,
      b => LPM_q_ivl_27418,
      c => LPM_d0_ivl_27426
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4267
  U4173: xnor_HPC2
    port map (
      a => LPM_q_ivl_27430,
      b => LPM_q_ivl_27437,
      c => LPM_d0_ivl_27445
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4268
  U4174: xnor_HPC2
    port map (
      a => LPM_q_ivl_27449,
      b => LPM_q_ivl_27456,
      c => LPM_d0_ivl_27468
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3110
  U4175: xor_HPC2
    port map (
      a => LPM_q_ivl_4853,
      b => LPM_q_ivl_4864,
      c => LPM_d0_ivl_4872
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3111
  U4176: xor_HPC2
    port map (
      a => LPM_q_ivl_4880,
      b => LPM_q_ivl_4891,
      c => LPM_d0_ivl_4899
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4269
  U4177: xor_HPC2
    port map (
      a => LPM_q_ivl_27472,
      b => LPM_q_ivl_27481,
      c => LPM_d0_ivl_27489
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4270
  U4178: xnor_HPC2
    port map (
      a => LPM_q_ivl_27495,
      b => LPM_q_ivl_27506,
      c => LPM_d0_ivl_27514
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4271
  U4179: xnor_HPC2
    port map (
      a => LPM_q_ivl_27518,
      b => LPM_q_ivl_27525,
      c => LPM_d0_ivl_27533
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4272
  U4180: xor_HPC2
    port map (
      a => LPM_q_ivl_27537,
      b => LPM_q_ivl_27546,
      c => LPM_d0_ivl_27554
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4273
  U4181: xnor_HPC2
    port map (
      a => LPM_q_ivl_27560,
      b => LPM_q_ivl_27571,
      c => LPM_d0_ivl_27579
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4274
  U4182: xnor_HPC2
    port map (
      a => LPM_q_ivl_27583,
      b => LPM_q_ivl_27590,
      c => LPM_d0_ivl_27598
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4275
  U4183: xnor_HPC2
    port map (
      a => LPM_q_ivl_27602,
      b => LPM_q_ivl_27609,
      c => LPM_d0_ivl_27617
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4276
  U4184: xnor_HPC2
    port map (
      a => LPM_q_ivl_27621,
      b => LPM_q_ivl_27628,
      c => LPM_d0_ivl_27640
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3112
  U4185: xor_HPC2
    port map (
      a => LPM_q_ivl_4907,
      b => LPM_q_ivl_4918,
      c => LPM_d0_ivl_4926
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4277
  U4186: xnor_HPC2
    port map (
      a => LPM_q_ivl_27644,
      b => LPM_q_ivl_27651,
      c => LPM_d0_ivl_27659
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4278
  U4187: xor_HPC2
    port map (
      a => LPM_q_ivl_27663,
      b => LPM_q_ivl_27672,
      c => LPM_d0_ivl_27680
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4279
  U4188: xor_HPC2
    port map (
      a => LPM_q_ivl_27686,
      b => LPM_q_ivl_27697,
      c => LPM_d0_ivl_27705
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4280
  U4189: xnor_HPC2
    port map (
      a => LPM_q_ivl_27709,
      b => LPM_q_ivl_27716,
      c => LPM_d0_ivl_27724
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4281
  U4190: xnor_HPC2
    port map (
      a => LPM_q_ivl_27728,
      b => LPM_q_ivl_27735,
      c => LPM_d0_ivl_27747
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3113
  U4191: xor_HPC2
    port map (
      a => LPM_q_ivl_4934,
      b => LPM_q_ivl_4945,
      c => LPM_d0_ivl_4953
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4282
  U4192: xnor_HPC2
    port map (
      a => LPM_q_ivl_27751,
      b => LPM_q_ivl_27758,
      c => LPM_d0_ivl_27766
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4283
  U4193: xor_HPC2
    port map (
      a => LPM_q_ivl_27770,
      b => LPM_q_ivl_27779,
      c => LPM_d0_ivl_27787
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4284
  U4194: xor_HPC2
    port map (
      a => LPM_q_ivl_27793,
      b => LPM_q_ivl_27804,
      c => LPM_d0_ivl_27812
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4285
  U4195: xnor_HPC2
    port map (
      a => LPM_q_ivl_27816,
      b => LPM_q_ivl_27823,
      c => LPM_d0_ivl_27831
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4286
  U4196: xnor_HPC2
    port map (
      a => LPM_q_ivl_27835,
      b => LPM_q_ivl_27842,
      c => LPM_d0_ivl_27854
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3114
  U4197: xor_HPC2
    port map (
      a => LPM_q_ivl_4961,
      b => LPM_q_ivl_4972,
      c => LPM_d0_ivl_4980
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4287
  U4198: xnor_HPC2
    port map (
      a => LPM_q_ivl_27858,
      b => LPM_q_ivl_27865,
      c => LPM_d0_ivl_27873
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4288
  U4199: xor_HPC2
    port map (
      a => LPM_q_ivl_27877,
      b => LPM_q_ivl_27886,
      c => LPM_d0_ivl_27894
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4289
  U4200: xnor_HPC2
    port map (
      a => LPM_q_ivl_27900,
      b => LPM_q_ivl_27911,
      c => LPM_d0_ivl_27919
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4290
  U4201: xnor_HPC2
    port map (
      a => LPM_q_ivl_27923,
      b => LPM_q_ivl_27930,
      c => LPM_d0_ivl_27938
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4291
  U4202: xnor_HPC2
    port map (
      a => LPM_q_ivl_27942,
      b => LPM_q_ivl_27949,
      c => LPM_d0_ivl_27961
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3115
  U4203: xor_HPC2
    port map (
      a => LPM_q_ivl_4988,
      b => LPM_q_ivl_4999,
      c => LPM_d0_ivl_5007
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4292
  U4204: xnor_HPC2
    port map (
      a => LPM_q_ivl_27965,
      b => LPM_q_ivl_27972,
      c => LPM_d0_ivl_27980
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4293
  U4205: xor_HPC2
    port map (
      a => LPM_q_ivl_27984,
      b => LPM_q_ivl_27993,
      c => LPM_d0_ivl_28001
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4294
  U4206: xnor_HPC2
    port map (
      a => LPM_q_ivl_28007,
      b => LPM_q_ivl_28018,
      c => LPM_d0_ivl_28026
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4295
  U4207: xnor_HPC2
    port map (
      a => LPM_q_ivl_28030,
      b => LPM_q_ivl_28037,
      c => LPM_d0_ivl_28045
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4296
  U4208: xnor_HPC2
    port map (
      a => LPM_q_ivl_28049,
      b => LPM_q_ivl_28056,
      c => LPM_d0_ivl_28068
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3116
  U4209: xor_HPC2
    port map (
      a => LPM_q_ivl_5015,
      b => LPM_q_ivl_5026,
      c => LPM_d0_ivl_5034
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4297
  U4210: xnor_HPC2
    port map (
      a => LPM_q_ivl_28072,
      b => LPM_q_ivl_28079,
      c => LPM_d0_ivl_28087
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4298
  U4211: xor_HPC2
    port map (
      a => LPM_q_ivl_28091,
      b => LPM_q_ivl_28100,
      c => LPM_d0_ivl_28108
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4299
  U4212: xor_HPC2
    port map (
      a => LPM_q_ivl_28114,
      b => LPM_q_ivl_28125,
      c => LPM_d0_ivl_28133
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4300
  U4213: xnor_HPC2
    port map (
      a => LPM_q_ivl_28137,
      b => LPM_q_ivl_28144,
      c => LPM_d0_ivl_28152
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4301
  U4214: xnor_HPC2
    port map (
      a => LPM_q_ivl_28156,
      b => LPM_q_ivl_28163,
      c => LPM_d0_ivl_28175
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3117
  U4215: xor_HPC2
    port map (
      a => LPM_q_ivl_5042,
      b => LPM_q_ivl_5053,
      c => LPM_d0_ivl_5061
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4302
  U4216: xnor_HPC2
    port map (
      a => LPM_q_ivl_28179,
      b => LPM_q_ivl_28186,
      c => LPM_d0_ivl_28194
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4303
  U4217: xor_HPC2
    port map (
      a => LPM_q_ivl_28198,
      b => LPM_q_ivl_28207,
      c => LPM_d0_ivl_28215
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4304
  U4218: xor_HPC2
    port map (
      a => LPM_q_ivl_28221,
      b => LPM_q_ivl_28232,
      c => LPM_d0_ivl_28240
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4305
  U4219: xnor_HPC2
    port map (
      a => LPM_q_ivl_28244,
      b => LPM_q_ivl_28251,
      c => LPM_d0_ivl_28259
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4306
  U4220: xnor_HPC2
    port map (
      a => LPM_q_ivl_28263,
      b => LPM_q_ivl_28270,
      c => LPM_d0_ivl_28282
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3118
  U4221: xor_HPC2
    port map (
      a => LPM_q_ivl_5069,
      b => LPM_q_ivl_5080,
      c => LPM_d0_ivl_5088
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4307
  U4222: xnor_HPC2
    port map (
      a => LPM_q_ivl_28286,
      b => LPM_q_ivl_28293,
      c => LPM_d0_ivl_28301
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4308
  U4223: xor_HPC2
    port map (
      a => LPM_q_ivl_28305,
      b => LPM_q_ivl_28314,
      c => LPM_d0_ivl_28322
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4309
  U4224: xnor_HPC2
    port map (
      a => LPM_q_ivl_28328,
      b => LPM_q_ivl_28339,
      c => LPM_d0_ivl_28347
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4310
  U4225: xnor_HPC2
    port map (
      a => LPM_q_ivl_28351,
      b => LPM_q_ivl_28358,
      c => LPM_d0_ivl_28366
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4311
  U4226: xnor_HPC2
    port map (
      a => LPM_q_ivl_28370,
      b => LPM_q_ivl_28377,
      c => LPM_d0_ivl_28389
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3119
  U4227: xor_HPC2
    port map (
      a => LPM_q_ivl_5096,
      b => LPM_q_ivl_5107,
      c => LPM_d0_ivl_5115
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4312
  U4228: xor_HPC2
    port map (
      a => LPM_q_ivl_28393,
      b => LPM_q_ivl_28402,
      c => LPM_d0_ivl_28410
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4313
  U4229: xnor_HPC2
    port map (
      a => LPM_q_ivl_28416,
      b => LPM_q_ivl_28427,
      c => LPM_d0_ivl_28435
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4314
  U4230: xnor_HPC2
    port map (
      a => LPM_q_ivl_28439,
      b => LPM_q_ivl_28446,
      c => LPM_d0_ivl_28454
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4315
  U4231: xnor_HPC2
    port map (
      a => LPM_q_ivl_28458,
      b => LPM_q_ivl_28465,
      c => LPM_d0_ivl_28473
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4316
  U4232: xnor_HPC2
    port map (
      a => LPM_q_ivl_28477,
      b => LPM_q_ivl_28484,
      c => LPM_d0_ivl_28496
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3120
  U4233: xor_HPC2
    port map (
      a => LPM_q_ivl_5123,
      b => LPM_q_ivl_5134,
      c => LPM_d0_ivl_5142
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4317
  U4234: xor_HPC2
    port map (
      a => LPM_q_ivl_28500,
      b => LPM_q_ivl_28509,
      c => LPM_d0_ivl_28517
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4318
  U4235: xnor_HPC2
    port map (
      a => LPM_q_ivl_28523,
      b => LPM_q_ivl_28534,
      c => LPM_d0_ivl_28542
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4319
  U4236: xnor_HPC2
    port map (
      a => LPM_q_ivl_28546,
      b => LPM_q_ivl_28553,
      c => LPM_d0_ivl_28561
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4320
  U4237: xnor_HPC2
    port map (
      a => LPM_q_ivl_28565,
      b => LPM_q_ivl_28572,
      c => LPM_d0_ivl_28580
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4321
  U4238: xnor_HPC2
    port map (
      a => LPM_q_ivl_28584,
      b => LPM_q_ivl_28591,
      c => LPM_d0_ivl_28603
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3121
  U4239: xor_HPC2
    port map (
      a => LPM_q_ivl_5150,
      b => LPM_q_ivl_5161,
      c => LPM_d0_ivl_5169
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4322
  U4240: xnor_HPC2
    port map (
      a => LPM_q_ivl_28607,
      b => LPM_q_ivl_28614,
      c => LPM_d0_ivl_28622
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4323
  U4241: xor_HPC2
    port map (
      a => LPM_q_ivl_28626,
      b => LPM_q_ivl_28635,
      c => LPM_d0_ivl_28643
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4324
  U4242: xnor_HPC2
    port map (
      a => LPM_q_ivl_28649,
      b => LPM_q_ivl_28660,
      c => LPM_d0_ivl_28668
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4325
  U4243: xnor_HPC2
    port map (
      a => LPM_q_ivl_28672,
      b => LPM_q_ivl_28679,
      c => LPM_d0_ivl_28687
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4326
  U4244: xnor_HPC2
    port map (
      a => LPM_q_ivl_28691,
      b => LPM_q_ivl_28698,
      c => LPM_d0_ivl_28710
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3122
  U4245: xor_HPC2
    port map (
      a => LPM_q_ivl_5177,
      b => LPM_q_ivl_5188,
      c => LPM_d0_ivl_5196
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4327
  U4246: xnor_HPC2
    port map (
      a => LPM_q_ivl_28714,
      b => LPM_q_ivl_28721,
      c => LPM_d0_ivl_28729
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4328
  U4247: xor_HPC2
    port map (
      a => LPM_q_ivl_28733,
      b => LPM_q_ivl_28742,
      c => LPM_d0_ivl_28750
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4329
  U4248: xnor_HPC2
    port map (
      a => LPM_q_ivl_28756,
      b => LPM_q_ivl_28767,
      c => LPM_d0_ivl_28775
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4330
  U4249: xnor_HPC2
    port map (
      a => LPM_q_ivl_28779,
      b => LPM_q_ivl_28786,
      c => LPM_d0_ivl_28794
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4331
  U4250: xnor_HPC2
    port map (
      a => LPM_q_ivl_28798,
      b => LPM_q_ivl_28805,
      c => LPM_d0_ivl_28817
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3123
  U4251: xor_HPC2
    port map (
      a => LPM_q_ivl_5204,
      b => LPM_q_ivl_5215,
      c => LPM_d0_ivl_5223
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4332
  U4252: xor_HPC2
    port map (
      a => LPM_q_ivl_28821,
      b => LPM_q_ivl_28830,
      c => LPM_d0_ivl_28838
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4333
  U4253: xnor_HPC2
    port map (
      a => LPM_q_ivl_28844,
      b => LPM_q_ivl_28855,
      c => LPM_d0_ivl_28863
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4334
  U4254: xnor_HPC2
    port map (
      a => LPM_q_ivl_28867,
      b => LPM_q_ivl_28874,
      c => LPM_d0_ivl_28882
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4335
  U4255: xnor_HPC2
    port map (
      a => LPM_q_ivl_28886,
      b => LPM_q_ivl_28893,
      c => LPM_d0_ivl_28901
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4336
  U4256: xnor_HPC2
    port map (
      a => LPM_q_ivl_28905,
      b => LPM_q_ivl_28912,
      c => LPM_d0_ivl_28924
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3124
  U4257: xor_HPC2
    port map (
      a => LPM_q_ivl_5231,
      b => LPM_q_ivl_5242,
      c => LPM_d0_ivl_5250
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4337
  U4258: xnor_HPC2
    port map (
      a => LPM_q_ivl_28928,
      b => LPM_q_ivl_28935,
      c => LPM_d0_ivl_28943
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4338
  U4259: xor_HPC2
    port map (
      a => LPM_q_ivl_28947,
      b => LPM_q_ivl_28956,
      c => LPM_d0_ivl_28964
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4339
  U4260: xor_HPC2
    port map (
      a => LPM_q_ivl_28970,
      b => LPM_q_ivl_28981,
      c => LPM_d0_ivl_28989
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4340
  U4261: xnor_HPC2
    port map (
      a => LPM_q_ivl_28993,
      b => LPM_q_ivl_29000,
      c => LPM_d0_ivl_29008
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4341
  U4262: xnor_HPC2
    port map (
      a => LPM_q_ivl_29012,
      b => LPM_q_ivl_29019,
      c => LPM_d0_ivl_29031
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3125
  U4263: xor_HPC2
    port map (
      a => LPM_q_ivl_5258,
      b => LPM_q_ivl_5269,
      c => LPM_d0_ivl_5277
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4342
  U4264: xor_HPC2
    port map (
      a => LPM_q_ivl_29035,
      b => LPM_q_ivl_29044,
      c => LPM_d0_ivl_29052
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4343
  U4265: xor_HPC2
    port map (
      a => LPM_q_ivl_29058,
      b => LPM_q_ivl_29069,
      c => LPM_d0_ivl_29077
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4344
  U4266: xnor_HPC2
    port map (
      a => LPM_q_ivl_29081,
      b => LPM_q_ivl_29088,
      c => LPM_d0_ivl_29096
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4345
  U4267: xor_HPC2
    port map (
      a => LPM_q_ivl_29100,
      b => LPM_q_ivl_29107,
      c => LPM_d0_ivl_29115
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4346
  U4268: xnor_HPC2
    port map (
      a => LPM_q_ivl_29119,
      b => LPM_q_ivl_29126,
      c => LPM_d0_ivl_29138
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3126
  U4269: xor_HPC2
    port map (
      a => LPM_q_ivl_5285,
      b => LPM_q_ivl_5296,
      c => LPM_d0_ivl_5304
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4347
  U4270: xor_HPC2
    port map (
      a => LPM_q_ivl_29142,
      b => LPM_q_ivl_29151,
      c => LPM_d0_ivl_29159
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4348
  U4271: xnor_HPC2
    port map (
      a => LPM_q_ivl_29165,
      b => LPM_q_ivl_29176,
      c => LPM_d0_ivl_29184
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4349
  U4272: xnor_HPC2
    port map (
      a => LPM_q_ivl_29188,
      b => LPM_q_ivl_29195,
      c => LPM_d0_ivl_29203
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4350
  U4273: xor_HPC2
    port map (
      a => LPM_q_ivl_29207,
      b => LPM_q_ivl_29214,
      c => LPM_d0_ivl_29222
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4351
  U4274: xnor_HPC2
    port map (
      a => LPM_q_ivl_29226,
      b => LPM_q_ivl_29233,
      c => LPM_d0_ivl_29245
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3127
  U4275: xor_HPC2
    port map (
      a => LPM_q_ivl_5312,
      b => LPM_q_ivl_5323,
      c => LPM_d0_ivl_5331
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4352
  U4276: xnor_HPC2
    port map (
      a => LPM_q_ivl_29249,
      b => LPM_q_ivl_29256,
      c => LPM_d0_ivl_29264
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4353
  U4277: xor_HPC2
    port map (
      a => LPM_q_ivl_29268,
      b => LPM_q_ivl_29277,
      c => LPM_d0_ivl_29285
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4354
  U4278: xor_HPC2
    port map (
      a => LPM_q_ivl_29291,
      b => LPM_q_ivl_29302,
      c => LPM_d0_ivl_29310
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4355
  U4279: xnor_HPC2
    port map (
      a => LPM_q_ivl_29314,
      b => LPM_q_ivl_29321,
      c => LPM_d0_ivl_29329
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4356
  U4280: xnor_HPC2
    port map (
      a => LPM_q_ivl_29333,
      b => LPM_q_ivl_29340,
      c => LPM_d0_ivl_29352
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3128
  U4281: xor_HPC2
    port map (
      a => LPM_q_ivl_5339,
      b => LPM_q_ivl_5350,
      c => LPM_d0_ivl_5358
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4357
  U4282: xnor_HPC2
    port map (
      a => LPM_q_ivl_29356,
      b => LPM_q_ivl_29363,
      c => LPM_d0_ivl_29371
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4358
  U4283: xor_HPC2
    port map (
      a => LPM_q_ivl_29375,
      b => LPM_q_ivl_29384,
      c => LPM_d0_ivl_29392
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4359
  U4284: xnor_HPC2
    port map (
      a => LPM_q_ivl_29398,
      b => LPM_q_ivl_29409,
      c => LPM_d0_ivl_29417
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4360
  U4285: xnor_HPC2
    port map (
      a => LPM_q_ivl_29421,
      b => LPM_q_ivl_29428,
      c => LPM_d0_ivl_29436
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4361
  U4286: xnor_HPC2
    port map (
      a => LPM_q_ivl_29440,
      b => LPM_q_ivl_29447,
      c => LPM_d0_ivl_29459
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3129
  U4287: xor_HPC2
    port map (
      a => LPM_q_ivl_5366,
      b => LPM_q_ivl_5377,
      c => LPM_d0_ivl_5385
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4362
  U4288: xor_HPC2
    port map (
      a => LPM_q_ivl_29463,
      b => LPM_q_ivl_29472,
      c => LPM_d0_ivl_29480
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4363
  U4289: xnor_HPC2
    port map (
      a => LPM_q_ivl_29486,
      b => LPM_q_ivl_29497,
      c => LPM_d0_ivl_29505
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4364
  U4290: xnor_HPC2
    port map (
      a => LPM_q_ivl_29509,
      b => LPM_q_ivl_29516,
      c => LPM_d0_ivl_29524
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4365
  U4291: xor_HPC2
    port map (
      a => LPM_q_ivl_29528,
      b => LPM_q_ivl_29535,
      c => LPM_d0_ivl_29543
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4366
  U4292: xnor_HPC2
    port map (
      a => LPM_q_ivl_29547,
      b => LPM_q_ivl_29554,
      c => LPM_d0_ivl_29566
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3130
  U4293: xor_HPC2
    port map (
      a => LPM_q_ivl_5393,
      b => LPM_q_ivl_5404,
      c => LPM_d0_ivl_5412
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4367
  U4294: xor_HPC2
    port map (
      a => LPM_q_ivl_29570,
      b => LPM_q_ivl_29579,
      c => LPM_d0_ivl_29587
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4368
  U4295: xnor_HPC2
    port map (
      a => LPM_q_ivl_29593,
      b => LPM_q_ivl_29604,
      c => LPM_d0_ivl_29612
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4369
  U4296: xnor_HPC2
    port map (
      a => LPM_q_ivl_29616,
      b => LPM_q_ivl_29623,
      c => LPM_d0_ivl_29631
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4370
  U4297: xor_HPC2
    port map (
      a => LPM_q_ivl_29635,
      b => LPM_q_ivl_29642,
      c => LPM_d0_ivl_29650
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4371
  U4298: xnor_HPC2
    port map (
      a => LPM_q_ivl_29654,
      b => LPM_q_ivl_29661,
      c => LPM_d0_ivl_29673
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3131
  U4299: xor_HPC2
    port map (
      a => LPM_q_ivl_5420,
      b => LPM_q_ivl_5431,
      c => LPM_d0_ivl_5439
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4372
  U4300: xnor_HPC2
    port map (
      a => LPM_q_ivl_29677,
      b => LPM_q_ivl_29684,
      c => LPM_d0_ivl_29692
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4373
  U4301: xor_HPC2
    port map (
      a => LPM_q_ivl_29696,
      b => LPM_q_ivl_29705,
      c => LPM_d0_ivl_29713
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4374
  U4302: xor_HPC2
    port map (
      a => LPM_q_ivl_29719,
      b => LPM_q_ivl_29730,
      c => LPM_d0_ivl_29738
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4375
  U4303: xnor_HPC2
    port map (
      a => LPM_q_ivl_29742,
      b => LPM_q_ivl_29749,
      c => LPM_d0_ivl_29757
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4376
  U4304: xnor_HPC2
    port map (
      a => LPM_q_ivl_29761,
      b => LPM_q_ivl_29768,
      c => LPM_d0_ivl_29780
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3132
  U4305: xor_HPC2
    port map (
      a => LPM_q_ivl_5447,
      b => LPM_q_ivl_5458,
      c => LPM_d0_ivl_5466
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4377
  U4306: xor_HPC2
    port map (
      a => LPM_q_ivl_29784,
      b => LPM_q_ivl_29793,
      c => LPM_d0_ivl_29801
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4378
  U4307: xor_HPC2
    port map (
      a => LPM_q_ivl_29807,
      b => LPM_q_ivl_29818,
      c => LPM_d0_ivl_29826
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4379
  U4308: xnor_HPC2
    port map (
      a => LPM_q_ivl_29830,
      b => LPM_q_ivl_29837,
      c => LPM_d0_ivl_29845
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4380
  U4309: xnor_HPC2
    port map (
      a => LPM_q_ivl_29849,
      b => LPM_q_ivl_29856,
      c => LPM_d0_ivl_29864
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4381
  U4310: xnor_HPC2
    port map (
      a => LPM_q_ivl_29868,
      b => LPM_q_ivl_29875,
      c => LPM_d0_ivl_29887
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3133
  U4311: xor_HPC2
    port map (
      a => LPM_q_ivl_5474,
      b => LPM_q_ivl_5485,
      c => LPM_d0_ivl_5493
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4382
  U4312: xor_HPC2
    port map (
      a => LPM_q_ivl_29891,
      b => LPM_q_ivl_29900,
      c => LPM_d0_ivl_29908
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4383
  U4313: xnor_HPC2
    port map (
      a => LPM_q_ivl_29914,
      b => LPM_q_ivl_29925,
      c => LPM_d0_ivl_29933
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4384
  U4314: xnor_HPC2
    port map (
      a => LPM_q_ivl_29937,
      b => LPM_q_ivl_29944,
      c => LPM_d0_ivl_29952
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4385
  U4315: xor_HPC2
    port map (
      a => LPM_q_ivl_29956,
      b => LPM_q_ivl_29963,
      c => LPM_d0_ivl_29971
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4386
  U4316: xnor_HPC2
    port map (
      a => LPM_q_ivl_29975,
      b => LPM_q_ivl_29982,
      c => LPM_d0_ivl_29994
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3134
  U4317: xor_HPC2
    port map (
      a => LPM_q_ivl_5501,
      b => LPM_q_ivl_5512,
      c => LPM_d0_ivl_5520
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4387
  U4318: xor_HPC2
    port map (
      a => LPM_q_ivl_29998,
      b => LPM_q_ivl_30007,
      c => LPM_d0_ivl_30015
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4388
  U4319: xnor_HPC2
    port map (
      a => LPM_q_ivl_30021,
      b => LPM_q_ivl_30032,
      c => LPM_d0_ivl_30040
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4389
  U4320: xnor_HPC2
    port map (
      a => LPM_q_ivl_30044,
      b => LPM_q_ivl_30051,
      c => LPM_d0_ivl_30059
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4390
  U4321: xnor_HPC2
    port map (
      a => LPM_q_ivl_30063,
      b => LPM_q_ivl_30070,
      c => LPM_d0_ivl_30078
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4391
  U4322: xnor_HPC2
    port map (
      a => LPM_q_ivl_30082,
      b => LPM_q_ivl_30089,
      c => LPM_d0_ivl_30101
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3135
  U4323: xor_HPC2
    port map (
      a => LPM_q_ivl_5528,
      b => LPM_q_ivl_5539,
      c => LPM_d0_ivl_5547
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4392
  U4324: xor_HPC2
    port map (
      a => LPM_q_ivl_30105,
      b => LPM_q_ivl_30114,
      c => LPM_d0_ivl_30122
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4393
  U4325: xnor_HPC2
    port map (
      a => LPM_q_ivl_30128,
      b => LPM_q_ivl_30139,
      c => LPM_d0_ivl_30147
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4394
  U4326: xnor_HPC2
    port map (
      a => LPM_q_ivl_30151,
      b => LPM_q_ivl_30158,
      c => LPM_d0_ivl_30166
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4395
  U4327: xnor_HPC2
    port map (
      a => LPM_q_ivl_30170,
      b => LPM_q_ivl_30177,
      c => LPM_d0_ivl_30185
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4396
  U4328: xnor_HPC2
    port map (
      a => LPM_q_ivl_30189,
      b => LPM_q_ivl_30196,
      c => LPM_d0_ivl_30208
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3136
  U4329: xor_HPC2
    port map (
      a => LPM_q_ivl_5555,
      b => LPM_q_ivl_5566,
      c => LPM_d0_ivl_5574
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4397
  U4330: xor_HPC2
    port map (
      a => LPM_q_ivl_30212,
      b => LPM_q_ivl_30221,
      c => LPM_d0_ivl_30229
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4398
  U4331: xor_HPC2
    port map (
      a => LPM_q_ivl_30235,
      b => LPM_q_ivl_30246,
      c => LPM_d0_ivl_30254
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4399
  U4332: xnor_HPC2
    port map (
      a => LPM_q_ivl_30258,
      b => LPM_q_ivl_30265,
      c => LPM_d0_ivl_30273
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4400
  U4333: xor_HPC2
    port map (
      a => LPM_q_ivl_30277,
      b => LPM_q_ivl_30284,
      c => LPM_d0_ivl_30292
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4401
  U4334: xnor_HPC2
    port map (
      a => LPM_q_ivl_30296,
      b => LPM_q_ivl_30303,
      c => LPM_d0_ivl_30315
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3137
  U4335: xor_HPC2
    port map (
      a => LPM_q_ivl_5582,
      b => LPM_q_ivl_5593,
      c => LPM_d0_ivl_5601
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4402
  U4336: xnor_HPC2
    port map (
      a => LPM_q_ivl_30321,
      b => LPM_q_ivl_30328,
      c => LPM_d0_ivl_30336
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4403
  U4337: xnor_HPC2
    port map (
      a => LPM_q_ivl_30344,
      b => LPM_q_ivl_30351,
      c => LPM_d0_ivl_30359
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4404
  U4338: xnor_HPC2
    port map (
      a => LPM_q_ivl_30363,
      b => LPM_q_ivl_30372,
      c => LPM_d0_ivl_30380
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4405
  U4339: xnor_HPC2
    port map (
      a => LPM_q_ivl_30384,
      b => LPM_q_ivl_30395,
      c => LPM_d0_ivl_30403
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4406
  U4340: xnor_HPC2
    port map (
      a => LPM_q_ivl_30407,
      b => LPM_q_ivl_30414,
      c => LPM_d0_ivl_30422
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4407
  U4341: xnor_HPC2
    port map (
      a => LPM_q_ivl_30426,
      b => LPM_q_ivl_30433,
      c => LPM_d0_ivl_30445
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4408
  U4342: xor_HPC2
    port map (
      a => LPM_q_ivl_30449,
      b => LPM_q_ivl_30456,
      c => LPM_d0_ivl_30464
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4409
  U4343: xnor_HPC2
    port map (
      a => LPM_q_ivl_30468,
      b => LPM_q_ivl_30475,
      c => LPM_d0_ivl_30487
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3138
  U4344: INV_X1
    port map (
      A => LPM_q_ivl_5602,
      ZN => n4068
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3139
  U4345: xnor_HPC2
    port map (
      a => LPM_q_ivl_5607,
      b => LPM_q_ivl_5616,
      c => LPM_d0_ivl_5626
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3140
  U4346: xor_HPC2
    port map (
      a => LPM_q_ivl_5634,
      b => LPM_q_ivl_5645,
      c => LPM_d0_ivl_5653
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4410
  U4347: xnor_HPC2
    port map (
      a => LPM_q_ivl_30491,
      b => LPM_q_ivl_30500,
      c => LPM_d0_ivl_30508
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4411
  U4348: xor_HPC2
    port map (
      a => LPM_q_ivl_30514,
      b => LPM_q_ivl_30525,
      c => LPM_d0_ivl_30533
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4412
  U4349: xnor_HPC2
    port map (
      a => LPM_q_ivl_30537,
      b => LPM_q_ivl_30544,
      c => LPM_d0_ivl_30552
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4413
  U4350: xnor_HPC2
    port map (
      a => LPM_q_ivl_30556,
      b => LPM_q_ivl_30563,
      c => LPM_d0_ivl_30571
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4414
  U4351: xnor_HPC2
    port map (
      a => LPM_q_ivl_30575,
      b => LPM_q_ivl_30582,
      c => LPM_d0_ivl_30594
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3141
  U4352: xor_HPC2
    port map (
      a => LPM_q_ivl_5661,
      b => LPM_q_ivl_5672,
      c => LPM_d0_ivl_5680
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4415
  U4353: xor_HPC2
    port map (
      a => LPM_q_ivl_30598,
      b => LPM_q_ivl_30607,
      c => LPM_d0_ivl_30615
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4416
  U4354: xnor_HPC2
    port map (
      a => LPM_q_ivl_30621,
      b => LPM_q_ivl_30632,
      c => LPM_d0_ivl_30640
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4417
  U4355: xnor_HPC2
    port map (
      a => LPM_q_ivl_30644,
      b => LPM_q_ivl_30651,
      c => LPM_d0_ivl_30659
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4418
  U4356: xnor_HPC2
    port map (
      a => LPM_q_ivl_30663,
      b => LPM_q_ivl_30670,
      c => LPM_d0_ivl_30678
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4419
  U4357: xnor_HPC2
    port map (
      a => LPM_q_ivl_30682,
      b => LPM_q_ivl_30689,
      c => LPM_d0_ivl_30701
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3142
  U4358: xor_HPC2
    port map (
      a => LPM_q_ivl_5688,
      b => LPM_q_ivl_5699,
      c => LPM_d0_ivl_5707
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4420
  U4359: xor_HPC2
    port map (
      a => LPM_q_ivl_30705,
      b => LPM_q_ivl_30714,
      c => LPM_d0_ivl_30722
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4421
  U4360: xnor_HPC2
    port map (
      a => LPM_q_ivl_30726,
      b => LPM_q_ivl_30735,
      c => LPM_d0_ivl_30743
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4422
  U4361: xnor_HPC2
    port map (
      a => LPM_q_ivl_30747,
      b => LPM_q_ivl_30758,
      c => LPM_d0_ivl_30766
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4423
  U4362: xnor_HPC2
    port map (
      a => LPM_q_ivl_30770,
      b => LPM_q_ivl_30777,
      c => LPM_d0_ivl_30785
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4424
  U4363: xnor_HPC2
    port map (
      a => LPM_q_ivl_30789,
      b => LPM_q_ivl_30796,
      c => LPM_d0_ivl_30808
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4425
  U4364: xor_HPC2
    port map (
      a => LPM_q_ivl_30812,
      b => LPM_q_ivl_30819,
      c => LPM_d0_ivl_30827
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4426
  U4365: xnor_HPC2
    port map (
      a => LPM_q_ivl_30831,
      b => LPM_q_ivl_30838,
      c => LPM_d0_ivl_30850
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3143
  U4366: xor_HPC2
    port map (
      a => LPM_q_ivl_5715,
      b => LPM_q_ivl_5726,
      c => LPM_d0_ivl_5734
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3144
  U4367: xnor_HPC2
    port map (
      a => LPM_q_ivl_5742,
      b => LPM_q_ivl_5749,
      c => LPM_d0_ivl_5757
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3145
  U4368: xor_HPC2
    port map (
      a => LPM_q_ivl_5765,
      b => LPM_q_ivl_5776,
      c => LPM_d0_ivl_5784
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4427
  U4369: xor_HPC2
    port map (
      a => LPM_q_ivl_30856,
      b => LPM_q_ivl_30863,
      c => LPM_d0_ivl_30871
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4428
  U4370: xor_HPC2
    port map (
      a => LPM_q_ivl_30875,
      b => LPM_q_ivl_30884,
      c => LPM_d0_ivl_30892
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4429
  U4371: xor_HPC2
    port map (
      a => LPM_q_ivl_30896,
      b => LPM_q_ivl_30903,
      c => LPM_d0_ivl_30911
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4430
  U4372: xnor_HPC2
    port map (
      a => LPM_q_ivl_30915,
      b => LPM_q_ivl_30922,
      c => LPM_d0_ivl_30934
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4431
  U4373: xnor_HPC2
    port map (
      a => LPM_q_ivl_30938,
      b => LPM_q_ivl_30945,
      c => LPM_d0_ivl_30953
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4432
  U4374: xnor_HPC2
    port map (
      a => LPM_q_ivl_30959,
      b => LPM_q_ivl_30970,
      c => LPM_d0_ivl_30978
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4433
  U4375: xnor_HPC2
    port map (
      a => LPM_q_ivl_30982,
      b => LPM_q_ivl_30989,
      c => LPM_d0_ivl_30997
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4434
  U4376: xnor_HPC2
    port map (
      a => LPM_q_ivl_31001,
      b => LPM_q_ivl_31008,
      c => LPM_d0_ivl_31020
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4435
  U4377: xor_HPC2
    port map (
      a => LPM_q_ivl_31024,
      b => LPM_q_ivl_31031,
      c => LPM_d0_ivl_31039
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4436
  U4378: xnor_HPC2
    port map (
      a => LPM_q_ivl_31043,
      b => LPM_q_ivl_31050,
      c => LPM_d0_ivl_31062
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3146
  U4379: INV_X1
    port map (
      A => LPM_q_ivl_5785,
      ZN => n4067
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3147
  U4380: XNOR2_X1
    port map (
      A => LPM_q_ivl_5787,
      B => n4067,
      ZN => n4206
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3148
  U4381: xor_HPC2
    port map (
      a => LPM_q_ivl_5796,
      b => LPM_q_ivl_5807,
      c => LPM_d0_ivl_5815
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4437
  U4382: xnor_HPC2
    port map (
      a => LPM_q_ivl_31068,
      b => LPM_q_ivl_31075,
      c => LPM_d0_ivl_31083
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4438
  U4383: xnor_HPC2
    port map (
      a => LPM_q_ivl_31089,
      b => LPM_q_ivl_31096,
      c => LPM_d0_ivl_31104
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4439
  U4384: xor_HPC2
    port map (
      a => LPM_q_ivl_31108,
      b => LPM_q_ivl_31117,
      c => LPM_d0_ivl_31125
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4440
  U4385: xnor_HPC2
    port map (
      a => LPM_q_ivl_31133,
      b => LPM_q_ivl_31140,
      c => LPM_d0_ivl_31148
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4441
  U4386: xnor_HPC2
    port map (
      a => LPM_q_ivl_31152,
      b => LPM_q_ivl_31159,
      c => LPM_d0_ivl_31167
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4442
  U4387: xnor_HPC2
    port map (
      a => LPM_q_ivl_31171,
      b => LPM_q_ivl_31178,
      c => LPM_d0_ivl_31190
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4443
  U4388: xnor_HPC2
    port map (
      a => LPM_q_ivl_31194,
      b => LPM_q_ivl_31201,
      c => LPM_d0_ivl_31209
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4444
  U4389: xnor_HPC2
    port map (
      a => LPM_q_ivl_31213,
      b => LPM_q_ivl_31220,
      c => LPM_d0_ivl_31232
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4445
  U4390: xor_HPC2
    port map (
      a => LPM_q_ivl_31236,
      b => LPM_q_ivl_31243,
      c => LPM_d0_ivl_31251
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4446
  U4391: xnor_HPC2
    port map (
      a => LPM_q_ivl_31255,
      b => LPM_q_ivl_31262,
      c => LPM_d0_ivl_31274
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3149
  U4392: xor_HPC2
    port map (
      a => LPM_q_ivl_5821,
      b => LPM_q_ivl_5828,
      c => LPM_d0_ivl_5838
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3150
  U4393: xnor_HPC2
    port map (
      a => LPM_q_ivl_5846,
      b => LPM_q_ivl_5857,
      c => LPM_d0_ivl_5865
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3151
  U4394: NAND2_X1
    port map (
      A1 => n4068,
      A2 => n4067,
      ZN => n4079
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3152
  U4395: XNOR2_X1
    port map (
      A => LPM_q_ivl_5866,
      B => n4079,
      ZN => n4087
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3153
  U4396: xnor_HPC2
    port map (
      a => LPM_q_ivl_5871,
      b => LPM_q_ivl_5880,
      c => LPM_d0_ivl_5888
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4447
  U4397: xnor_HPC2
    port map (
      a => LPM_q_ivl_31280,
      b => LPM_q_ivl_31287,
      c => LPM_d0_ivl_31295
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4448
  U4398: xnor_HPC2
    port map (
      a => LPM_q_ivl_31301,
      b => LPM_q_ivl_31312,
      c => LPM_d0_ivl_31320
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4449
  U4399: xnor_HPC2
    port map (
      a => LPM_q_ivl_31324,
      b => LPM_q_ivl_31331,
      c => LPM_d0_ivl_31339
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4450
  U4400: xnor_HPC2
    port map (
      a => LPM_q_ivl_31343,
      b => LPM_q_ivl_31350,
      c => LPM_d0_ivl_31358
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4451
  U4401: xnor_HPC2
    port map (
      a => LPM_q_ivl_31362,
      b => LPM_q_ivl_31369,
      c => LPM_d0_ivl_31381
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4452
  U4402: xnor_HPC2
    port map (
      a => LPM_q_ivl_31385,
      b => LPM_q_ivl_31392,
      c => LPM_d0_ivl_31400
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4453
  U4403: xnor_HPC2
    port map (
      a => LPM_q_ivl_31404,
      b => LPM_q_ivl_31411,
      c => LPM_d0_ivl_31423
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4454
  U4404: xnor_HPC2
    port map (
      a => LPM_q_ivl_31427,
      b => LPM_q_ivl_31434,
      c => LPM_d0_ivl_31442
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4455
  U4405: xnor_HPC2
    port map (
      a => LPM_q_ivl_31446,
      b => LPM_q_ivl_31453,
      c => LPM_d0_ivl_31465
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3154
  U4406: NAND2_X1
    port map (
      A1 => LPM_q_ivl_5889,
      A2 => n4079,
      ZN => n4080
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3155
  U4407: XNOR2_X1
    port map (
      A => LPM_q_ivl_5891,
      B => n4080,
      ZN => n4084
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3156
  U4408: xor_HPC2
    port map (
      a => LPM_q_ivl_5898,
      b => LPM_q_ivl_5909,
      c => LPM_d0_ivl_5917
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3157
  U4409: xnor_HPC2
    port map (
      a => LPM_q_ivl_5925,
      b => LPM_q_ivl_5932,
      c => LPM_d0_ivl_5940
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4456
  U4410: xnor_HPC2
    port map (
      a => LPM_q_ivl_31471,
      b => LPM_q_ivl_31478,
      c => LPM_d0_ivl_31486
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4457
  U4411: xnor_HPC2
    port map (
      a => LPM_q_ivl_31490,
      b => LPM_q_ivl_31497,
      c => LPM_d0_ivl_31505
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4458
  U4412: xnor_HPC2
    port map (
      a => LPM_q_ivl_31509,
      b => LPM_q_ivl_31516,
      c => LPM_d0_ivl_31528
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4459
  U4413: xnor_HPC2
    port map (
      a => LPM_q_ivl_31532,
      b => LPM_q_ivl_31539,
      c => LPM_d0_ivl_31547
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4460
  U4414: xnor_HPC2
    port map (
      a => LPM_q_ivl_31551,
      b => LPM_q_ivl_31558,
      c => LPM_d0_ivl_31570
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3158
  U4415: xnor_HPC2
    port map (
      a => LPM_q_ivl_5946,
      b => LPM_q_ivl_5957,
      c => LPM_d0_ivl_5965
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3159
  U4416: xnor_HPC2
    port map (
      a => LPM_q_ivl_5969,
      b => LPM_q_ivl_5980,
      c => LPM_d0_ivl_5988
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3160
  U4417: xor_HPC2
    port map (
      a => LPM_q_ivl_5996,
      b => LPM_q_ivl_6007,
      c => LPM_d0_ivl_6015
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3161
  U4418: xnor_HPC2
    port map (
      a => LPM_q_ivl_6021,
      b => LPM_q_ivl_6028,
      c => LPM_d0_ivl_6036
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4461
  U4419: xor_HPC2
    port map (
      a => LPM_q_ivl_31574,
      b => LPM_q_ivl_31583,
      c => LPM_d0_ivl_31591
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4462
  U4420: xnor_HPC2
    port map (
      a => LPM_q_ivl_31595,
      b => LPM_q_ivl_31602,
      c => LPM_d0_ivl_31610
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4463
  U4421: xnor_HPC2
    port map (
      a => LPM_q_ivl_31614,
      b => LPM_q_ivl_31623,
      c => LPM_d0_ivl_31631
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4464
  U4422: xnor_HPC2
    port map (
      a => LPM_q_ivl_31635,
      b => LPM_q_ivl_31642,
      c => LPM_d0_ivl_31654
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4465
  U4423: xnor_HPC2
    port map (
      a => LPM_q_ivl_31660,
      b => LPM_q_ivl_31671,
      c => LPM_d0_ivl_31679
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4466
  U4424: xnor_HPC2
    port map (
      a => LPM_q_ivl_31683,
      b => LPM_q_ivl_31690,
      c => LPM_d0_ivl_31698
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4467
  U4425: xnor_HPC2
    port map (
      a => LPM_q_ivl_31702,
      b => LPM_q_ivl_31709,
      c => LPM_d0_ivl_31717
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4468
  U4426: xnor_HPC2
    port map (
      a => LPM_q_ivl_31721,
      b => LPM_q_ivl_31728,
      c => LPM_d0_ivl_31740
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4469
  U4427: xnor_HPC2
    port map (
      a => LPM_q_ivl_31744,
      b => LPM_q_ivl_31751,
      c => LPM_d0_ivl_31759
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4470
  U4428: xnor_HPC2
    port map (
      a => LPM_q_ivl_31763,
      b => LPM_q_ivl_31770,
      c => LPM_d0_ivl_31782
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4471
  U4429: xnor_HPC2
    port map (
      a => LPM_q_ivl_31786,
      b => LPM_q_ivl_31793,
      c => LPM_d0_ivl_31801
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4472
  U4430: xnor_HPC2
    port map (
      a => LPM_q_ivl_31805,
      b => LPM_q_ivl_31812,
      c => LPM_d0_ivl_31824
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4473
  U4431: xnor_HPC2
    port map (
      a => LPM_q_ivl_31828,
      b => LPM_q_ivl_31835,
      c => LPM_d0_ivl_31843
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3162
  U4432: xnor_HPC2
    port map (
      a => LPM_q_ivl_6044,
      b => LPM_q_ivl_6055,
      c => LPM_d0_ivl_6063
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4474
  U4433: xnor_HPC2
    port map (
      a => LPM_q_ivl_31849,
      b => LPM_q_ivl_31856,
      c => LPM_d0_ivl_31864
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4475
  U4434: xnor_HPC2
    port map (
      a => LPM_q_ivl_31872,
      b => LPM_q_ivl_31879,
      c => LPM_d0_ivl_31887
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4476
  U4435: xnor_HPC2
    port map (
      a => LPM_q_ivl_31891,
      b => LPM_q_ivl_31898,
      c => LPM_d0_ivl_31910
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4477
  U4436: xor_HPC2
    port map (
      a => LPM_q_ivl_31914,
      b => LPM_q_ivl_31921,
      c => LPM_d0_ivl_31929
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4478
  U4437: xnor_HPC2
    port map (
      a => LPM_q_ivl_31933,
      b => LPM_q_ivl_31940,
      c => LPM_d0_ivl_31948
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4479
  U4438: xnor_HPC2
    port map (
      a => LPM_q_ivl_31956,
      b => LPM_q_ivl_31963,
      c => LPM_d0_ivl_31975
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:3163
  U4439: xor_HPC2
    port map (
      a => LPM_q_ivl_6069,
      b => LPM_q_ivl_6076,
      c => LPM_d0_ivl_6084
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4480
  U4440: xor_HPC2
    port map (
      a => LPM_q_ivl_31979,
      b => LPM_q_ivl_31986,
      c => LPM_d0_ivl_31994
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4481
  U4441: xnor_HPC2
    port map (
      a => LPM_q_ivl_31998,
      b => LPM_q_ivl_32005,
      c => LPM_d0_ivl_32017
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4482
  U4442: xor_HPC2
    port map (
      a => LPM_q_ivl_32021,
      b => LPM_q_ivl_32028,
      c => LPM_d0_ivl_32036
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4483
  U4443: xnor_HPC2
    port map (
      a => LPM_q_ivl_32040,
      b => LPM_q_ivl_32047,
      c => LPM_d0_ivl_32059
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4484
  U4444: xor_HPC2
    port map (
      a => LPM_q_ivl_32063,
      b => LPM_q_ivl_32070,
      c => LPM_d0_ivl_32078
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4485
  U4445: xnor_HPC2
    port map (
      a => LPM_q_ivl_32082,
      b => LPM_q_ivl_32089,
      c => LPM_d0_ivl_32101
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4486
  U4446: xor_HPC2
    port map (
      a => LPM_q_ivl_32105,
      b => LPM_q_ivl_32112,
      c => LPM_d0_ivl_32120
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4487
  U4447: xnor_HPC2
    port map (
      a => LPM_q_ivl_32124,
      b => LPM_q_ivl_32131,
      c => LPM_d0_ivl_32143
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4488
  U4448: xor_HPC2
    port map (
      a => LPM_q_ivl_32147,
      b => LPM_q_ivl_32154,
      c => LPM_d0_ivl_32162
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4489
  U4449: xnor_HPC2
    port map (
      a => LPM_q_ivl_32166,
      b => LPM_q_ivl_32173,
      c => LPM_d0_ivl_32185
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4490
  U4450: xor_HPC2
    port map (
      a => LPM_q_ivl_32189,
      b => LPM_q_ivl_32196,
      c => LPM_d0_ivl_32204
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4491
  U4451: xnor_HPC2
    port map (
      a => LPM_q_ivl_32208,
      b => LPM_q_ivl_32215,
      c => LPM_d0_ivl_32227
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4492
  U4452: xor_HPC2
    port map (
      a => LPM_q_ivl_32231,
      b => LPM_q_ivl_32238,
      c => LPM_d0_ivl_32246
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4493
  U4453: xnor_HPC2
    port map (
      a => LPM_q_ivl_32250,
      b => LPM_q_ivl_32257,
      c => LPM_d0_ivl_32269
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4494
  U4454: xor_HPC2
    port map (
      a => LPM_q_ivl_32273,
      b => LPM_q_ivl_32280,
      c => LPM_d0_ivl_32288
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4495
  U4455: xnor_HPC2
    port map (
      a => LPM_q_ivl_32292,
      b => LPM_q_ivl_32299,
      c => LPM_d0_ivl_32311
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4496
  U4456: xor_HPC2
    port map (
      a => LPM_q_ivl_32315,
      b => LPM_q_ivl_32322,
      c => LPM_d0_ivl_32330
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4497
  U4457: xnor_HPC2
    port map (
      a => LPM_q_ivl_32334,
      b => LPM_q_ivl_32341,
      c => LPM_d0_ivl_32353
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4498
  U4458: xor_HPC2
    port map (
      a => LPM_q_ivl_32357,
      b => LPM_q_ivl_32364,
      c => LPM_d0_ivl_32372
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4499
  U4459: xnor_HPC2
    port map (
      a => LPM_q_ivl_32376,
      b => LPM_q_ivl_32383,
      c => LPM_d0_ivl_32395
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4500
  U4460: xor_HPC2
    port map (
      a => LPM_q_ivl_32399,
      b => LPM_q_ivl_32406,
      c => LPM_d0_ivl_32414
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4501
  U4461: xnor_HPC2
    port map (
      a => LPM_q_ivl_32418,
      b => LPM_q_ivl_32425,
      c => LPM_d0_ivl_32437
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4502
  U4462: xor_HPC2
    port map (
      a => LPM_q_ivl_32441,
      b => LPM_q_ivl_32448,
      c => LPM_d0_ivl_32456
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4503
  U4463: xnor_HPC2
    port map (
      a => LPM_q_ivl_32460,
      b => LPM_q_ivl_32467,
      c => LPM_d0_ivl_32479
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4504
  U4464: xor_HPC2
    port map (
      a => LPM_q_ivl_32483,
      b => LPM_q_ivl_32490,
      c => LPM_d0_ivl_32498
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4505
  U4465: xnor_HPC2
    port map (
      a => LPM_q_ivl_32502,
      b => LPM_q_ivl_32509,
      c => LPM_d0_ivl_32521
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4506
  U4466: xor_HPC2
    port map (
      a => LPM_q_ivl_32525,
      b => LPM_q_ivl_32532,
      c => LPM_d0_ivl_32540
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4507
  U4467: xnor_HPC2
    port map (
      a => LPM_q_ivl_32544,
      b => LPM_q_ivl_32551,
      c => LPM_d0_ivl_32563
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4508
  U4468: xor_HPC2
    port map (
      a => LPM_q_ivl_32567,
      b => LPM_q_ivl_32574,
      c => LPM_d0_ivl_32582
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4509
  U4469: xnor_HPC2
    port map (
      a => LPM_q_ivl_32586,
      b => LPM_q_ivl_32593,
      c => LPM_d0_ivl_32605
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4510
  U4470: xor_HPC2
    port map (
      a => LPM_q_ivl_32609,
      b => LPM_q_ivl_32616,
      c => LPM_d0_ivl_32624
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4511
  U4471: xnor_HPC2
    port map (
      a => LPM_q_ivl_32628,
      b => LPM_q_ivl_32635,
      c => LPM_d0_ivl_32647
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4512
  U4472: xor_HPC2
    port map (
      a => LPM_q_ivl_32651,
      b => LPM_q_ivl_32658,
      c => LPM_d0_ivl_32666
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4513
  U4473: xnor_HPC2
    port map (
      a => LPM_q_ivl_32670,
      b => LPM_q_ivl_32677,
      c => LPM_d0_ivl_32689
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4514
  U4474: xor_HPC2
    port map (
      a => LPM_q_ivl_32693,
      b => LPM_q_ivl_32700,
      c => LPM_d0_ivl_32708
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4515
  U4475: xnor_HPC2
    port map (
      a => LPM_q_ivl_32712,
      b => LPM_q_ivl_32719,
      c => LPM_d0_ivl_32731
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4516
  U4476: xor_HPC2
    port map (
      a => LPM_q_ivl_32735,
      b => LPM_q_ivl_32742,
      c => LPM_d0_ivl_32750
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4517
  U4477: xnor_HPC2
    port map (
      a => LPM_q_ivl_32754,
      b => LPM_q_ivl_32761,
      c => LPM_d0_ivl_32773
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4518
  U4478: xor_HPC2
    port map (
      a => LPM_q_ivl_32777,
      b => LPM_q_ivl_32784,
      c => LPM_d0_ivl_32792
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4519
  U4479: xnor_HPC2
    port map (
      a => LPM_q_ivl_32796,
      b => LPM_q_ivl_32803,
      c => LPM_d0_ivl_32815
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4520
  U4480: xor_HPC2
    port map (
      a => LPM_q_ivl_32819,
      b => LPM_q_ivl_32826,
      c => LPM_d0_ivl_32834
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4521
  U4481: xnor_HPC2
    port map (
      a => LPM_q_ivl_32838,
      b => LPM_q_ivl_32845,
      c => LPM_d0_ivl_32857
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4522
  U4482: xor_HPC2
    port map (
      a => LPM_q_ivl_32861,
      b => LPM_q_ivl_32868,
      c => LPM_d0_ivl_32876
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4523
  U4483: xnor_HPC2
    port map (
      a => LPM_q_ivl_32880,
      b => LPM_q_ivl_32887,
      c => LPM_d0_ivl_32899
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4524
  U4484: xor_HPC2
    port map (
      a => LPM_q_ivl_32903,
      b => LPM_q_ivl_32910,
      c => LPM_d0_ivl_32918
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4525
  U4485: xnor_HPC2
    port map (
      a => LPM_q_ivl_32922,
      b => LPM_q_ivl_32929,
      c => LPM_d0_ivl_32941
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4526
  U4486: xor_HPC2
    port map (
      a => LPM_q_ivl_32945,
      b => LPM_q_ivl_32952,
      c => LPM_d0_ivl_32960
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4527
  U4487: xnor_HPC2
    port map (
      a => LPM_q_ivl_32964,
      b => LPM_q_ivl_32971,
      c => LPM_d0_ivl_32983
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4528
  U4488: xor_HPC2
    port map (
      a => LPM_q_ivl_32987,
      b => LPM_q_ivl_32994,
      c => LPM_d0_ivl_33002
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4529
  U4489: xnor_HPC2
    port map (
      a => LPM_q_ivl_33006,
      b => LPM_q_ivl_33013,
      c => LPM_d0_ivl_33025
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4530
  U4490: xor_HPC2
    port map (
      a => LPM_q_ivl_33029,
      b => LPM_q_ivl_33036,
      c => LPM_d0_ivl_33044
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4531
  U4491: xnor_HPC2
    port map (
      a => LPM_q_ivl_33048,
      b => LPM_q_ivl_33055,
      c => LPM_d0_ivl_33067
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4532
  U4492: xor_HPC2
    port map (
      a => LPM_q_ivl_33071,
      b => LPM_q_ivl_33078,
      c => LPM_d0_ivl_33086
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4533
  U4493: xnor_HPC2
    port map (
      a => LPM_q_ivl_33090,
      b => LPM_q_ivl_33097,
      c => LPM_d0_ivl_33109
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4534
  U4494: xor_HPC2
    port map (
      a => LPM_q_ivl_33113,
      b => LPM_q_ivl_33120,
      c => LPM_d0_ivl_33128
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4535
  U4495: xnor_HPC2
    port map (
      a => LPM_q_ivl_33132,
      b => LPM_q_ivl_33139,
      c => LPM_d0_ivl_33151
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4536
  U4496: xor_HPC2
    port map (
      a => LPM_q_ivl_33155,
      b => LPM_q_ivl_33162,
      c => LPM_d0_ivl_33170
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4537
  U4497: xnor_HPC2
    port map (
      a => LPM_q_ivl_33174,
      b => LPM_q_ivl_33181,
      c => LPM_d0_ivl_33193
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4538
  U4498: xor_HPC2
    port map (
      a => LPM_q_ivl_33197,
      b => LPM_q_ivl_33204,
      c => LPM_d0_ivl_33212
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4539
  U4499: xnor_HPC2
    port map (
      a => LPM_q_ivl_33216,
      b => LPM_q_ivl_33223,
      c => LPM_d0_ivl_33235
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4540
  U4500: xor_HPC2
    port map (
      a => LPM_q_ivl_33239,
      b => LPM_q_ivl_33246,
      c => LPM_d0_ivl_33254
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4541
  U4501: xnor_HPC2
    port map (
      a => LPM_q_ivl_33258,
      b => LPM_q_ivl_33265,
      c => LPM_d0_ivl_33277
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4542
  U4502: xor_HPC2
    port map (
      a => LPM_q_ivl_33281,
      b => LPM_q_ivl_33288,
      c => LPM_d0_ivl_33296
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4543
  U4503: xnor_HPC2
    port map (
      a => LPM_q_ivl_33300,
      b => LPM_q_ivl_33307,
      c => LPM_d0_ivl_33319
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4544
  U4504: xor_HPC2
    port map (
      a => LPM_q_ivl_33323,
      b => LPM_q_ivl_33330,
      c => LPM_d0_ivl_33338
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4545
  U4505: xnor_HPC2
    port map (
      a => LPM_q_ivl_33342,
      b => LPM_q_ivl_33349,
      c => LPM_d0_ivl_33361
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4546
  U4506: xor_HPC2
    port map (
      a => LPM_q_ivl_33365,
      b => LPM_q_ivl_33372,
      c => LPM_d0_ivl_33380
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4547
  U4507: xnor_HPC2
    port map (
      a => LPM_q_ivl_33384,
      b => LPM_q_ivl_33391,
      c => LPM_d0_ivl_33403
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4548
  U4508: xor_HPC2
    port map (
      a => LPM_q_ivl_33407,
      b => LPM_q_ivl_33414,
      c => LPM_d0_ivl_33422
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4549
  U4509: xnor_HPC2
    port map (
      a => LPM_q_ivl_33426,
      b => LPM_q_ivl_33433,
      c => LPM_d0_ivl_33445
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4550
  U4510: xor_HPC2
    port map (
      a => LPM_q_ivl_33449,
      b => LPM_q_ivl_33456,
      c => LPM_d0_ivl_33464
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4551
  U4511: xnor_HPC2
    port map (
      a => LPM_q_ivl_33468,
      b => LPM_q_ivl_33475,
      c => LPM_d0_ivl_33487
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4552
  U4512: xor_HPC2
    port map (
      a => LPM_q_ivl_33491,
      b => LPM_q_ivl_33498,
      c => LPM_d0_ivl_33506
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4553
  U4513: xnor_HPC2
    port map (
      a => LPM_q_ivl_33510,
      b => LPM_q_ivl_33517,
      c => LPM_d0_ivl_33529
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4554
  U4514: xor_HPC2
    port map (
      a => LPM_q_ivl_33533,
      b => LPM_q_ivl_33540,
      c => LPM_d0_ivl_33548
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4555
  U4515: xnor_HPC2
    port map (
      a => LPM_q_ivl_33552,
      b => LPM_q_ivl_33559,
      c => LPM_d0_ivl_33571
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4556
  U4516: xor_HPC2
    port map (
      a => LPM_q_ivl_33575,
      b => LPM_q_ivl_33582,
      c => LPM_d0_ivl_33590
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4557
  U4517: xnor_HPC2
    port map (
      a => LPM_q_ivl_33594,
      b => LPM_q_ivl_33601,
      c => LPM_d0_ivl_33613
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4558
  U4518: xor_HPC2
    port map (
      a => LPM_q_ivl_33617,
      b => LPM_q_ivl_33624,
      c => LPM_d0_ivl_33632
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4559
  U4519: xnor_HPC2
    port map (
      a => LPM_q_ivl_33636,
      b => LPM_q_ivl_33643,
      c => LPM_d0_ivl_33655
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4560
  U4520: xor_HPC2
    port map (
      a => LPM_q_ivl_33659,
      b => LPM_q_ivl_33666,
      c => LPM_d0_ivl_33674
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4561
  U4521: xnor_HPC2
    port map (
      a => LPM_q_ivl_33678,
      b => LPM_q_ivl_33685,
      c => LPM_d0_ivl_33697
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4562
  U4522: xor_HPC2
    port map (
      a => LPM_q_ivl_33701,
      b => LPM_q_ivl_33708,
      c => LPM_d0_ivl_33716
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4563
  U4523: xnor_HPC2
    port map (
      a => LPM_q_ivl_33720,
      b => LPM_q_ivl_33727,
      c => LPM_d0_ivl_33739
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4564
  U4524: xor_HPC2
    port map (
      a => LPM_q_ivl_33743,
      b => LPM_q_ivl_33750,
      c => LPM_d0_ivl_33758
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4565
  U4525: xnor_HPC2
    port map (
      a => LPM_q_ivl_33762,
      b => LPM_q_ivl_33769,
      c => LPM_d0_ivl_33781
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4566
  U4526: xor_HPC2
    port map (
      a => LPM_q_ivl_33785,
      b => LPM_q_ivl_33792,
      c => LPM_d0_ivl_33800
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4567
  U4527: xnor_HPC2
    port map (
      a => LPM_q_ivl_33804,
      b => LPM_q_ivl_33811,
      c => LPM_d0_ivl_33823
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4568
  U4528: xor_HPC2
    port map (
      a => LPM_q_ivl_33827,
      b => LPM_q_ivl_33834,
      c => LPM_d0_ivl_33842
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4569
  U4529: xnor_HPC2
    port map (
      a => LPM_q_ivl_33846,
      b => LPM_q_ivl_33853,
      c => LPM_d0_ivl_33865
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4570
  U4530: xor_HPC2
    port map (
      a => LPM_q_ivl_33869,
      b => LPM_q_ivl_33876,
      c => LPM_d0_ivl_33884
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4571
  U4531: xnor_HPC2
    port map (
      a => LPM_q_ivl_33888,
      b => LPM_q_ivl_33895,
      c => LPM_d0_ivl_33907
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4572
  U4532: xor_HPC2
    port map (
      a => LPM_q_ivl_33911,
      b => LPM_q_ivl_33918,
      c => LPM_d0_ivl_33926
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4573
  U4533: xnor_HPC2
    port map (
      a => LPM_q_ivl_33930,
      b => LPM_q_ivl_33937,
      c => LPM_d0_ivl_33949
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4574
  U4534: xor_HPC2
    port map (
      a => LPM_q_ivl_33953,
      b => LPM_q_ivl_33960,
      c => LPM_d0_ivl_33968
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4575
  U4535: xnor_HPC2
    port map (
      a => LPM_q_ivl_33972,
      b => LPM_q_ivl_33979,
      c => LPM_d0_ivl_33991
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4576
  U4536: xor_HPC2
    port map (
      a => LPM_q_ivl_33995,
      b => LPM_q_ivl_34002,
      c => LPM_d0_ivl_34010
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4577
  U4537: xnor_HPC2
    port map (
      a => LPM_q_ivl_34014,
      b => LPM_q_ivl_34021,
      c => LPM_d0_ivl_34033
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4578
  U4538: xnor_HPC2
    port map (
      a => LPM_q_ivl_34037,
      b => LPM_q_ivl_34044,
      c => LPM_d0_ivl_34052
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4579
  U4539: xnor_HPC2
    port map (
      a => LPM_q_ivl_34056,
      b => LPM_q_ivl_34063,
      c => LPM_d0_ivl_34075
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4580
  U4540: xnor_HPC2
    port map (
      a => LPM_q_ivl_34079,
      b => LPM_q_ivl_34086,
      c => LPM_d0_ivl_34094
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4581
  U4541: xnor_HPC2
    port map (
      a => LPM_q_ivl_34098,
      b => LPM_q_ivl_34105,
      c => LPM_d0_ivl_34117
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4582
  U4542: xnor_HPC2
    port map (
      a => LPM_q_ivl_34121,
      b => LPM_q_ivl_34128,
      c => LPM_d0_ivl_34136
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4583
  U4543: xnor_HPC2
    port map (
      a => LPM_q_ivl_34142,
      b => LPM_q_ivl_34149,
      c => LPM_d0_ivl_34157
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4584
  U4544: xnor_HPC2
    port map (
      a => LPM_q_ivl_34161,
      b => LPM_q_ivl_34168,
      c => LPM_d0_ivl_34180
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4585
  U4545: xor_HPC2
    port map (
      a => LPM_q_ivl_34184,
      b => LPM_q_ivl_34193,
      c => LPM_d0_ivl_34201
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4586
  U4546: xnor_HPC2
    port map (
      a => LPM_q_ivl_34205,
      b => LPM_q_ivl_34212,
      c => LPM_d0_ivl_34220
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4587
  U4547: xnor_HPC2
    port map (
      a => LPM_q_ivl_34224,
      b => LPM_q_ivl_34231,
      c => LPM_d0_ivl_34243
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4588
  U4548: xnor_HPC2
    port map (
      a => LPM_q_ivl_34247,
      b => LPM_q_ivl_34254,
      c => LPM_d0_ivl_34262
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4589
  U4549: xnor_HPC2
    port map (
      a => LPM_q_ivl_34266,
      b => LPM_q_ivl_34273,
      c => LPM_d0_ivl_34285
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4590
  U4550: xnor_HPC2
    port map (
      a => LPM_q_ivl_34289,
      b => LPM_q_ivl_34296,
      c => LPM_d0_ivl_34304
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4591
  U4551: xnor_HPC2
    port map (
      a => LPM_q_ivl_34308,
      b => LPM_q_ivl_34315,
      c => LPM_d0_ivl_34327
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4592
  U4552: xnor_HPC2
    port map (
      a => LPM_q_ivl_34331,
      b => LPM_q_ivl_34338,
      c => LPM_d0_ivl_34346
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4593
  U4553: xnor_HPC2
    port map (
      a => LPM_q_ivl_34350,
      b => LPM_q_ivl_34357,
      c => LPM_d0_ivl_34369
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4594
  U4554: xor_HPC2
    port map (
      a => LPM_q_ivl_34373,
      b => LPM_q_ivl_34380,
      c => LPM_d0_ivl_34388
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4595
  U4555: xnor_HPC2
    port map (
      a => LPM_q_ivl_34392,
      b => LPM_q_ivl_34399,
      c => LPM_d0_ivl_34411
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4596
  U4556: xor_HPC2
    port map (
      a => LPM_q_ivl_34415,
      b => LPM_q_ivl_34422,
      c => LPM_d0_ivl_34430
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4597
  U4557: xnor_HPC2
    port map (
      a => LPM_q_ivl_34434,
      b => LPM_q_ivl_34441,
      c => LPM_d0_ivl_34453
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4598
  U4558: xor_HPC2
    port map (
      a => LPM_q_ivl_34459,
      b => LPM_q_ivl_34470,
      c => LPM_d0_ivl_34478
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4599
  U4559: xnor_HPC2
    port map (
      a => LPM_q_ivl_34482,
      b => LPM_q_ivl_34489,
      c => LPM_d0_ivl_34497
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4600
  U4560: xnor_HPC2
    port map (
      a => LPM_q_ivl_34501,
      b => LPM_q_ivl_34508,
      c => LPM_d0_ivl_34516
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4601
  U4561: xnor_HPC2
    port map (
      a => LPM_q_ivl_34520,
      b => LPM_q_ivl_34527,
      c => LPM_d0_ivl_34539
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4602
  U4562: xnor_HPC2
    port map (
      a => LPM_q_ivl_34543,
      b => LPM_q_ivl_34550,
      c => LPM_d0_ivl_34558
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4603
  U4563: xnor_HPC2
    port map (
      a => LPM_q_ivl_34562,
      b => LPM_q_ivl_34569,
      c => LPM_d0_ivl_34581
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4604
  U4564: xnor_HPC2
    port map (
      a => LPM_q_ivl_34585,
      b => LPM_q_ivl_34592,
      c => LPM_d0_ivl_34600
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4605
  U4565: xnor_HPC2
    port map (
      a => LPM_q_ivl_34604,
      b => LPM_q_ivl_34611,
      c => LPM_d0_ivl_34623
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4606
  U4566: xnor_HPC2
    port map (
      a => LPM_q_ivl_34629,
      b => LPM_q_ivl_34640,
      c => LPM_d0_ivl_34648
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4607
  U4567: xnor_HPC2
    port map (
      a => LPM_q_ivl_34652,
      b => LPM_q_ivl_34659,
      c => LPM_d0_ivl_34667
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4608
  U4568: xnor_HPC2
    port map (
      a => LPM_q_ivl_34671,
      b => LPM_q_ivl_34678,
      c => LPM_d0_ivl_34686
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4609
  U4569: xnor_HPC2
    port map (
      a => LPM_q_ivl_34690,
      b => LPM_q_ivl_34697,
      c => LPM_d0_ivl_34709
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4610
  U4570: xnor_HPC2
    port map (
      a => LPM_q_ivl_34713,
      b => LPM_q_ivl_34720,
      c => LPM_d0_ivl_34728
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4611
  U4571: xnor_HPC2
    port map (
      a => LPM_q_ivl_34732,
      b => LPM_q_ivl_34739,
      c => LPM_d0_ivl_34751
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4612
  U4572: xnor_HPC2
    port map (
      a => LPM_q_ivl_34755,
      b => LPM_q_ivl_34762,
      c => LPM_d0_ivl_34770
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4613
  U4573: xnor_HPC2
    port map (
      a => LPM_q_ivl_34774,
      b => LPM_q_ivl_34781,
      c => LPM_d0_ivl_34793
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4614
  U4574: xor_HPC2
    port map (
      a => LPM_q_ivl_34799,
      b => LPM_q_ivl_34810,
      c => LPM_d0_ivl_34818
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4615
  U4575: xnor_HPC2
    port map (
      a => LPM_q_ivl_34822,
      b => LPM_q_ivl_34829,
      c => LPM_d0_ivl_34837
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4616
  U4576: xnor_HPC2
    port map (
      a => LPM_q_ivl_34841,
      b => LPM_q_ivl_34848,
      c => LPM_d0_ivl_34856
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4617
  U4577: xnor_HPC2
    port map (
      a => LPM_q_ivl_34860,
      b => LPM_q_ivl_34867,
      c => LPM_d0_ivl_34879
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4618
  U4578: xor_HPC2
    port map (
      a => LPM_q_ivl_34883,
      b => LPM_q_ivl_34890,
      c => LPM_d0_ivl_34898
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4619
  U4579: xnor_HPC2
    port map (
      a => LPM_q_ivl_34902,
      b => LPM_q_ivl_34909,
      c => LPM_d0_ivl_34921
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4620
  U4580: xor_HPC2
    port map (
      a => LPM_q_ivl_34925,
      b => LPM_q_ivl_34932,
      c => LPM_d0_ivl_34940
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4621
  U4581: xnor_HPC2
    port map (
      a => LPM_q_ivl_34944,
      b => LPM_q_ivl_34951,
      c => LPM_d0_ivl_34963
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4622
  U4582: xnor_HPC2
    port map (
      a => LPM_q_ivl_34969,
      b => LPM_q_ivl_34980,
      c => LPM_d0_ivl_34988
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4623
  U4583: xnor_HPC2
    port map (
      a => LPM_q_ivl_34992,
      b => LPM_q_ivl_34999,
      c => LPM_d0_ivl_35007
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4624
  U4584: xnor_HPC2
    port map (
      a => LPM_q_ivl_35011,
      b => LPM_q_ivl_35018,
      c => LPM_d0_ivl_35026
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4625
  U4585: xnor_HPC2
    port map (
      a => LPM_q_ivl_35030,
      b => LPM_q_ivl_35037,
      c => LPM_d0_ivl_35049
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4626
  U4586: xnor_HPC2
    port map (
      a => LPM_q_ivl_35053,
      b => LPM_q_ivl_35060,
      c => LPM_d0_ivl_35068
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4627
  U4587: xnor_HPC2
    port map (
      a => LPM_q_ivl_35072,
      b => LPM_q_ivl_35079,
      c => LPM_d0_ivl_35091
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4628
  U4588: xnor_HPC2
    port map (
      a => LPM_q_ivl_35095,
      b => LPM_q_ivl_35102,
      c => LPM_d0_ivl_35110
    );
  
  -- Generated from instantiation at Ascon/Ascon128v12_first_order/src_rtl/Asconp_HPC2_ClockGating_d1.v:4629
  U4589: xnor_HPC2
    port map (
      a => LPM_q_ivl_35114,
      b => LPM_q_ivl_35121,
      c => LPM_d0_ivl_35133
    );
  tmp_ivl_10048 <= '0';
  tmp_ivl_10055 <= '0';
  tmp_ivl_1006 <= '0';
  tmp_ivl_10071 <= '0';
  tmp_ivl_10080 <= '0';
  tmp_ivl_10096 <= '0';
  tmp_ivl_10103 <= '0';
  tmp_ivl_10115 <= '0';
  tmp_ivl_10122 <= '0';
  tmp_ivl_10140 <= '0';
  tmp_ivl_10151 <= '0';
  tmp_ivl_10165 <= '0';
  tmp_ivl_10172 <= '0';
  tmp_ivl_10184 <= '0';
  tmp_ivl_10191 <= '0';
  tmp_ivl_10205 <= '0';
  tmp_ivl_10216 <= '0';
  tmp_ivl_10230 <= '0';
  tmp_ivl_1024 <= '0';
  tmp_ivl_10241 <= '0';
  tmp_ivl_10257 <= '0';
  tmp_ivl_10264 <= '0';
  tmp_ivl_10276 <= '0';
  tmp_ivl_10283 <= '0';
  tmp_ivl_10295 <= '0';
  tmp_ivl_10302 <= '0';
  tmp_ivl_10316 <= '0';
  tmp_ivl_10327 <= '0';
  tmp_ivl_10341 <= '0';
  tmp_ivl_1035 <= '0';
  tmp_ivl_10352 <= '0';
  tmp_ivl_10368 <= '0';
  tmp_ivl_10375 <= '0';
  tmp_ivl_10387 <= '0';
  tmp_ivl_10394 <= '0';
  tmp_ivl_10406 <= '0';
  tmp_ivl_10413 <= '0';
  tmp_ivl_10431 <= '0';
  tmp_ivl_10442 <= '0';
  tmp_ivl_10456 <= '0';
  tmp_ivl_10463 <= '0';
  tmp_ivl_10475 <= '0';
  tmp_ivl_10482 <= '0';
  tmp_ivl_10496 <= '0';
  tmp_ivl_10507 <= '0';
  tmp_ivl_10521 <= '0';
  tmp_ivl_1053 <= '0';
  tmp_ivl_10532 <= '0';
  tmp_ivl_10548 <= '0';
  tmp_ivl_10555 <= '0';
  tmp_ivl_10567 <= '0';
  tmp_ivl_10574 <= '0';
  tmp_ivl_10586 <= '0';
  tmp_ivl_10593 <= '0';
  tmp_ivl_10607 <= '0';
  tmp_ivl_10618 <= '0';
  tmp_ivl_10632 <= '0';
  tmp_ivl_1064 <= '0';
  tmp_ivl_10643 <= '0';
  tmp_ivl_10659 <= '0';
  tmp_ivl_10666 <= '0';
  tmp_ivl_10678 <= '0';
  tmp_ivl_10685 <= '0';
  tmp_ivl_10697 <= '0';
  tmp_ivl_107 <= '0';
  tmp_ivl_10704 <= '0';
  tmp_ivl_10720 <= '0';
  tmp_ivl_10727 <= '0';
  tmp_ivl_10743 <= '0';
  tmp_ivl_10752 <= '0';
  tmp_ivl_10768 <= '0';
  tmp_ivl_10775 <= '0';
  tmp_ivl_10787 <= '0';
  tmp_ivl_10794 <= '0';
  tmp_ivl_10810 <= '0';
  tmp_ivl_10817 <= '0';
  tmp_ivl_1082 <= '0';
  tmp_ivl_10833 <= '0';
  tmp_ivl_10842 <= '0';
  tmp_ivl_10858 <= '0';
  tmp_ivl_10865 <= '0';
  tmp_ivl_10877 <= '0';
  tmp_ivl_10884 <= '0';
  tmp_ivl_10904 <= '0';
  tmp_ivl_10913 <= '0';
  tmp_ivl_10929 <= '0';
  tmp_ivl_1093 <= '0';
  tmp_ivl_10936 <= '0';
  tmp_ivl_10948 <= '0';
  tmp_ivl_10955 <= '0';
  tmp_ivl_10971 <= '0';
  tmp_ivl_10980 <= '0';
  tmp_ivl_10996 <= '0';
  tmp_ivl_11003 <= '0';
  tmp_ivl_11015 <= '0';
  tmp_ivl_11022 <= '0';
  tmp_ivl_11040 <= '0';
  tmp_ivl_11051 <= '0';
  tmp_ivl_11065 <= '0';
  tmp_ivl_11076 <= '0';
  tmp_ivl_11092 <= '0';
  tmp_ivl_11099 <= '0';
  tmp_ivl_1111 <= '0';
  tmp_ivl_11111 <= '0';
  tmp_ivl_11118 <= '0';
  tmp_ivl_11132 <= '0';
  tmp_ivl_11143 <= '0';
  tmp_ivl_11157 <= '0';
  tmp_ivl_11164 <= '0';
  tmp_ivl_11176 <= '0';
  tmp_ivl_11183 <= '0';
  tmp_ivl_11195 <= '0';
  tmp_ivl_11202 <= '0';
  tmp_ivl_11216 <= '0';
  tmp_ivl_1122 <= '0';
  tmp_ivl_11227 <= '0';
  tmp_ivl_11241 <= '0';
  tmp_ivl_11252 <= '0';
  tmp_ivl_11268 <= '0';
  tmp_ivl_11275 <= '0';
  tmp_ivl_11287 <= '0';
  tmp_ivl_11294 <= '0';
  tmp_ivl_11306 <= '0';
  tmp_ivl_11313 <= '0';
  tmp_ivl_11331 <= '0';
  tmp_ivl_11342 <= '0';
  tmp_ivl_11356 <= '0';
  tmp_ivl_11367 <= '0';
  tmp_ivl_11383 <= '0';
  tmp_ivl_11390 <= '0';
  tmp_ivl_1140 <= '0';
  tmp_ivl_11402 <= '0';
  tmp_ivl_11409 <= '0';
  tmp_ivl_11421 <= '0';
  tmp_ivl_11428 <= '0';
  tmp_ivl_11442 <= '0';
  tmp_ivl_11453 <= '0';
  tmp_ivl_11467 <= '0';
  tmp_ivl_11474 <= '0';
  tmp_ivl_11486 <= '0';
  tmp_ivl_11493 <= '0';
  tmp_ivl_11505 <= '0';
  tmp_ivl_1151 <= '0';
  tmp_ivl_11512 <= '0';
  tmp_ivl_11530 <= '0';
  tmp_ivl_11541 <= '0';
  tmp_ivl_11555 <= '0';
  tmp_ivl_11566 <= '0';
  tmp_ivl_11582 <= '0';
  tmp_ivl_11589 <= '0';
  tmp_ivl_11601 <= '0';
  tmp_ivl_11608 <= '0';
  tmp_ivl_11620 <= '0';
  tmp_ivl_11627 <= '0';
  tmp_ivl_11641 <= '0';
  tmp_ivl_11652 <= '0';
  tmp_ivl_11666 <= '0';
  tmp_ivl_11677 <= '0';
  tmp_ivl_1169 <= '0';
  tmp_ivl_11693 <= '0';
  tmp_ivl_11700 <= '0';
  tmp_ivl_11712 <= '0';
  tmp_ivl_11719 <= '0';
  tmp_ivl_11731 <= '0';
  tmp_ivl_11738 <= '0';
  tmp_ivl_11754 <= '0';
  tmp_ivl_11761 <= '0';
  tmp_ivl_11777 <= '0';
  tmp_ivl_11786 <= '0';
  tmp_ivl_1180 <= '0';
  tmp_ivl_11802 <= '0';
  tmp_ivl_11809 <= '0';
  tmp_ivl_11821 <= '0';
  tmp_ivl_11828 <= '0';
  tmp_ivl_11844 <= '0';
  tmp_ivl_11851 <= '0';
  tmp_ivl_11863 <= '0';
  tmp_ivl_11870 <= '0';
  tmp_ivl_11888 <= '0';
  tmp_ivl_11899 <= '0';
  tmp_ivl_11913 <= '0';
  tmp_ivl_11924 <= '0';
  tmp_ivl_11940 <= '0';
  tmp_ivl_11947 <= '0';
  tmp_ivl_11959 <= '0';
  tmp_ivl_11966 <= '0';
  tmp_ivl_11978 <= '0';
  tmp_ivl_1198 <= '0';
  tmp_ivl_11985 <= '0';
  tmp_ivl_11999 <= '0';
  tmp_ivl_12010 <= '0';
  tmp_ivl_12024 <= '0';
  tmp_ivl_12031 <= '0';
  tmp_ivl_12043 <= '0';
  tmp_ivl_12050 <= '0';
  tmp_ivl_12062 <= '0';
  tmp_ivl_12069 <= '0';
  tmp_ivl_12085 <= '0';
  tmp_ivl_1209 <= '0';
  tmp_ivl_12092 <= '0';
  tmp_ivl_12108 <= '0';
  tmp_ivl_12117 <= '0';
  tmp_ivl_12133 <= '0';
  tmp_ivl_12140 <= '0';
  tmp_ivl_12152 <= '0';
  tmp_ivl_12159 <= '0';
  tmp_ivl_12177 <= '0';
  tmp_ivl_12188 <= '0';
  tmp_ivl_12200 <= '0';
  tmp_ivl_12207 <= '0';
  tmp_ivl_12221 <= '0';
  tmp_ivl_12232 <= '0';
  tmp_ivl_12244 <= '0';
  tmp_ivl_12251 <= '0';
  tmp_ivl_12263 <= '0';
  tmp_ivl_1227 <= '0';
  tmp_ivl_12270 <= '0';
  tmp_ivl_12282 <= '0';
  tmp_ivl_12289 <= '0';
  tmp_ivl_12301 <= '0';
  tmp_ivl_12308 <= '0';
  tmp_ivl_12328 <= '0';
  tmp_ivl_12337 <= '0';
  tmp_ivl_12353 <= '0';
  tmp_ivl_12360 <= '0';
  tmp_ivl_12372 <= '0';
  tmp_ivl_12379 <= '0';
  tmp_ivl_1238 <= '0';
  tmp_ivl_12395 <= '0';
  tmp_ivl_12404 <= '0';
  tmp_ivl_12420 <= '0';
  tmp_ivl_12427 <= '0';
  tmp_ivl_12439 <= '0';
  tmp_ivl_12446 <= '0';
  tmp_ivl_12462 <= '0';
  tmp_ivl_12469 <= '0';
  tmp_ivl_12481 <= '0';
  tmp_ivl_12488 <= '0';
  tmp_ivl_125 <= '0';
  tmp_ivl_12504 <= '0';
  tmp_ivl_12511 <= '0';
  tmp_ivl_12527 <= '0';
  tmp_ivl_12536 <= '0';
  tmp_ivl_12552 <= '0';
  tmp_ivl_12559 <= '0';
  tmp_ivl_1256 <= '0';
  tmp_ivl_12571 <= '0';
  tmp_ivl_12578 <= '0';
  tmp_ivl_12596 <= '0';
  tmp_ivl_12607 <= '0';
  tmp_ivl_12621 <= '0';
  tmp_ivl_12632 <= '0';
  tmp_ivl_12648 <= '0';
  tmp_ivl_12655 <= '0';
  tmp_ivl_12667 <= '0';
  tmp_ivl_1267 <= '0';
  tmp_ivl_12674 <= '0';
  tmp_ivl_12686 <= '0';
  tmp_ivl_12693 <= '0';
  tmp_ivl_12707 <= '0';
  tmp_ivl_12718 <= '0';
  tmp_ivl_12732 <= '0';
  tmp_ivl_12743 <= '0';
  tmp_ivl_12759 <= '0';
  tmp_ivl_12766 <= '0';
  tmp_ivl_12778 <= '0';
  tmp_ivl_12785 <= '0';
  tmp_ivl_12797 <= '0';
  tmp_ivl_12804 <= '0';
  tmp_ivl_12822 <= '0';
  tmp_ivl_12833 <= '0';
  tmp_ivl_12847 <= '0';
  tmp_ivl_1285 <= '0';
  tmp_ivl_12854 <= '0';
  tmp_ivl_12866 <= '0';
  tmp_ivl_12873 <= '0';
  tmp_ivl_12887 <= '0';
  tmp_ivl_12894 <= '0';
  tmp_ivl_12906 <= '0';
  tmp_ivl_12913 <= '0';
  tmp_ivl_12925 <= '0';
  tmp_ivl_12932 <= '0';
  tmp_ivl_12946 <= '0';
  tmp_ivl_12957 <= '0';
  tmp_ivl_1296 <= '0';
  tmp_ivl_12971 <= '0';
  tmp_ivl_12982 <= '0';
  tmp_ivl_12998 <= '0';
  tmp_ivl_13005 <= '0';
  tmp_ivl_13017 <= '0';
  tmp_ivl_13024 <= '0';
  tmp_ivl_13036 <= '0';
  tmp_ivl_13043 <= '0';
  tmp_ivl_13059 <= '0';
  tmp_ivl_13066 <= '0';
  tmp_ivl_13082 <= '0';
  tmp_ivl_13091 <= '0';
  tmp_ivl_13107 <= '0';
  tmp_ivl_13114 <= '0';
  tmp_ivl_13126 <= '0';
  tmp_ivl_13133 <= '0';
  tmp_ivl_1314 <= '0';
  tmp_ivl_13149 <= '0';
  tmp_ivl_13156 <= '0';
  tmp_ivl_13172 <= '0';
  tmp_ivl_13181 <= '0';
  tmp_ivl_13197 <= '0';
  tmp_ivl_13204 <= '0';
  tmp_ivl_13216 <= '0';
  tmp_ivl_13223 <= '0';
  tmp_ivl_13239 <= '0';
  tmp_ivl_13246 <= '0';
  tmp_ivl_1325 <= '0';
  tmp_ivl_13258 <= '0';
  tmp_ivl_13265 <= '0';
  tmp_ivl_13283 <= '0';
  tmp_ivl_13294 <= '0';
  tmp_ivl_13308 <= '0';
  tmp_ivl_13319 <= '0';
  tmp_ivl_13335 <= '0';
  tmp_ivl_13342 <= '0';
  tmp_ivl_13354 <= '0';
  tmp_ivl_13361 <= '0';
  tmp_ivl_13373 <= '0';
  tmp_ivl_13380 <= '0';
  tmp_ivl_13394 <= '0';
  tmp_ivl_13405 <= '0';
  tmp_ivl_13419 <= '0';
  tmp_ivl_1343 <= '0';
  tmp_ivl_13430 <= '0';
  tmp_ivl_13446 <= '0';
  tmp_ivl_13453 <= '0';
  tmp_ivl_13465 <= '0';
  tmp_ivl_13472 <= '0';
  tmp_ivl_13484 <= '0';
  tmp_ivl_13491 <= '0';
  tmp_ivl_13509 <= '0';
  tmp_ivl_13520 <= '0';
  tmp_ivl_13534 <= '0';
  tmp_ivl_1354 <= '0';
  tmp_ivl_13545 <= '0';
  tmp_ivl_13561 <= '0';
  tmp_ivl_13568 <= '0';
  tmp_ivl_13580 <= '0';
  tmp_ivl_13587 <= '0';
  tmp_ivl_136 <= '0';
  tmp_ivl_13601 <= '0';
  tmp_ivl_13612 <= '0';
  tmp_ivl_13626 <= '0';
  tmp_ivl_13633 <= '0';
  tmp_ivl_13645 <= '0';
  tmp_ivl_13652 <= '0';
  tmp_ivl_13664 <= '0';
  tmp_ivl_13671 <= '0';
  tmp_ivl_13685 <= '0';
  tmp_ivl_13696 <= '0';
  tmp_ivl_13710 <= '0';
  tmp_ivl_13717 <= '0';
  tmp_ivl_1372 <= '0';
  tmp_ivl_13729 <= '0';
  tmp_ivl_13736 <= '0';
  tmp_ivl_13748 <= '0';
  tmp_ivl_13755 <= '0';
  tmp_ivl_13771 <= '0';
  tmp_ivl_13778 <= '0';
  tmp_ivl_13794 <= '0';
  tmp_ivl_13803 <= '0';
  tmp_ivl_13819 <= '0';
  tmp_ivl_13826 <= '0';
  tmp_ivl_1383 <= '0';
  tmp_ivl_13838 <= '0';
  tmp_ivl_13845 <= '0';
  tmp_ivl_13861 <= '0';
  tmp_ivl_13868 <= '0';
  tmp_ivl_13880 <= '0';
  tmp_ivl_13887 <= '0';
  tmp_ivl_13903 <= '0';
  tmp_ivl_13910 <= '0';
  tmp_ivl_13922 <= '0';
  tmp_ivl_13929 <= '0';
  tmp_ivl_13943 <= '0';
  tmp_ivl_13954 <= '0';
  tmp_ivl_13966 <= '0';
  tmp_ivl_13973 <= '0';
  tmp_ivl_13985 <= '0';
  tmp_ivl_13992 <= '0';
  tmp_ivl_1401 <= '0';
  tmp_ivl_14010 <= '0';
  tmp_ivl_14021 <= '0';
  tmp_ivl_14037 <= '0';
  tmp_ivl_14044 <= '0';
  tmp_ivl_14056 <= '0';
  tmp_ivl_14063 <= '0';
  tmp_ivl_14075 <= '0';
  tmp_ivl_14082 <= '0';
  tmp_ivl_14096 <= '0';
  tmp_ivl_14107 <= '0';
  tmp_ivl_1412 <= '0';
  tmp_ivl_14121 <= '0';
  tmp_ivl_14132 <= '0';
  tmp_ivl_14148 <= '0';
  tmp_ivl_14155 <= '0';
  tmp_ivl_14167 <= '0';
  tmp_ivl_14174 <= '0';
  tmp_ivl_14186 <= '0';
  tmp_ivl_14193 <= '0';
  tmp_ivl_14211 <= '0';
  tmp_ivl_14222 <= '0';
  tmp_ivl_14234 <= '0';
  tmp_ivl_14241 <= '0';
  tmp_ivl_14255 <= '0';
  tmp_ivl_14266 <= '0';
  tmp_ivl_14278 <= '0';
  tmp_ivl_14285 <= '0';
  tmp_ivl_14297 <= '0';
  tmp_ivl_1430 <= '0';
  tmp_ivl_14304 <= '0';
  tmp_ivl_14316 <= '0';
  tmp_ivl_14323 <= '0';
  tmp_ivl_14335 <= '0';
  tmp_ivl_14342 <= '0';
  tmp_ivl_14360 <= '0';
  tmp_ivl_14371 <= '0';
  tmp_ivl_14387 <= '0';
  tmp_ivl_14394 <= '0';
  tmp_ivl_14406 <= '0';
  tmp_ivl_1441 <= '0';
  tmp_ivl_14413 <= '0';
  tmp_ivl_14425 <= '0';
  tmp_ivl_14432 <= '0';
  tmp_ivl_14446 <= '0';
  tmp_ivl_14457 <= '0';
  tmp_ivl_14473 <= '0';
  tmp_ivl_14480 <= '0';
  tmp_ivl_14492 <= '0';
  tmp_ivl_14499 <= '0';
  tmp_ivl_14511 <= '0';
  tmp_ivl_14518 <= '0';
  tmp_ivl_14534 <= '0';
  tmp_ivl_14541 <= '0';
  tmp_ivl_14553 <= '0';
  tmp_ivl_14560 <= '0';
  tmp_ivl_14578 <= '0';
  tmp_ivl_14589 <= '0';
  tmp_ivl_1459 <= '0';
  tmp_ivl_14605 <= '0';
  tmp_ivl_14614 <= '0';
  tmp_ivl_14626 <= '0';
  tmp_ivl_14633 <= '0';
  tmp_ivl_14647 <= '0';
  tmp_ivl_14658 <= '0';
  tmp_ivl_14670 <= '0';
  tmp_ivl_14677 <= '0';
  tmp_ivl_14689 <= '0';
  tmp_ivl_14696 <= '0';
  tmp_ivl_1470 <= '0';
  tmp_ivl_14708 <= '0';
  tmp_ivl_14715 <= '0';
  tmp_ivl_14727 <= '0';
  tmp_ivl_14734 <= '0';
  tmp_ivl_14750 <= '0';
  tmp_ivl_14757 <= '0';
  tmp_ivl_14773 <= '0';
  tmp_ivl_14780 <= '0';
  tmp_ivl_14792 <= '0';
  tmp_ivl_14799 <= '0';
  tmp_ivl_14817 <= '0';
  tmp_ivl_14828 <= '0';
  tmp_ivl_14842 <= '0';
  tmp_ivl_14853 <= '0';
  tmp_ivl_14869 <= '0';
  tmp_ivl_14876 <= '0';
  tmp_ivl_1488 <= '0';
  tmp_ivl_14888 <= '0';
  tmp_ivl_14895 <= '0';
  tmp_ivl_14909 <= '0';
  tmp_ivl_14920 <= '0';
  tmp_ivl_14936 <= '0';
  tmp_ivl_14943 <= '0';
  tmp_ivl_14955 <= '0';
  tmp_ivl_14962 <= '0';
  tmp_ivl_14974 <= '0';
  tmp_ivl_14981 <= '0';
  tmp_ivl_1499 <= '0';
  tmp_ivl_14995 <= '0';
  tmp_ivl_15006 <= '0';
  tmp_ivl_15020 <= '0';
  tmp_ivl_15027 <= '0';
  tmp_ivl_15039 <= '0';
  tmp_ivl_15046 <= '0';
  tmp_ivl_15058 <= '0';
  tmp_ivl_15065 <= '0';
  tmp_ivl_15081 <= '0';
  tmp_ivl_15088 <= '0';
  tmp_ivl_15100 <= '0';
  tmp_ivl_15107 <= '0';
  tmp_ivl_15123 <= '0';
  tmp_ivl_15130 <= '0';
  tmp_ivl_15142 <= '0';
  tmp_ivl_15149 <= '0';
  tmp_ivl_15167 <= '0';
  tmp_ivl_1517 <= '0';
  tmp_ivl_15178 <= '0';
  tmp_ivl_15190 <= '0';
  tmp_ivl_15197 <= '0';
  tmp_ivl_15209 <= '0';
  tmp_ivl_15216 <= '0';
  tmp_ivl_15228 <= '0';
  tmp_ivl_15235 <= '0';
  tmp_ivl_15247 <= '0';
  tmp_ivl_15254 <= '0';
  tmp_ivl_15266 <= '0';
  tmp_ivl_15273 <= '0';
  tmp_ivl_1528 <= '0';
  tmp_ivl_15291 <= '0';
  tmp_ivl_15302 <= '0';
  tmp_ivl_15318 <= '0';
  tmp_ivl_15325 <= '0';
  tmp_ivl_15337 <= '0';
  tmp_ivl_15344 <= '0';
  tmp_ivl_15356 <= '0';
  tmp_ivl_15363 <= '0';
  tmp_ivl_15377 <= '0';
  tmp_ivl_15384 <= '0';
  tmp_ivl_15396 <= '0';
  tmp_ivl_154 <= '0';
  tmp_ivl_15403 <= '0';
  tmp_ivl_15415 <= '0';
  tmp_ivl_15422 <= '0';
  tmp_ivl_15438 <= '0';
  tmp_ivl_15445 <= '0';
  tmp_ivl_15457 <= '0';
  tmp_ivl_1546 <= '0';
  tmp_ivl_15464 <= '0';
  tmp_ivl_15480 <= '0';
  tmp_ivl_15487 <= '0';
  tmp_ivl_15503 <= '0';
  tmp_ivl_15512 <= '0';
  tmp_ivl_15528 <= '0';
  tmp_ivl_15535 <= '0';
  tmp_ivl_15547 <= '0';
  tmp_ivl_15554 <= '0';
  tmp_ivl_1557 <= '0';
  tmp_ivl_15570 <= '0';
  tmp_ivl_15577 <= '0';
  tmp_ivl_15589 <= '0';
  tmp_ivl_15596 <= '0';
  tmp_ivl_15612 <= '0';
  tmp_ivl_15619 <= '0';
  tmp_ivl_15631 <= '0';
  tmp_ivl_15638 <= '0';
  tmp_ivl_15654 <= '0';
  tmp_ivl_15661 <= '0';
  tmp_ivl_15675 <= '0';
  tmp_ivl_15686 <= '0';
  tmp_ivl_15700 <= '0';
  tmp_ivl_15711 <= '0';
  tmp_ivl_15727 <= '0';
  tmp_ivl_15734 <= '0';
  tmp_ivl_15746 <= '0';
  tmp_ivl_1575 <= '0';
  tmp_ivl_15753 <= '0';
  tmp_ivl_15765 <= '0';
  tmp_ivl_15772 <= '0';
  tmp_ivl_15788 <= '0';
  tmp_ivl_15795 <= '0';
  tmp_ivl_15809 <= '0';
  tmp_ivl_15820 <= '0';
  tmp_ivl_15834 <= '0';
  tmp_ivl_15845 <= '0';
  tmp_ivl_1586 <= '0';
  tmp_ivl_15861 <= '0';
  tmp_ivl_15868 <= '0';
  tmp_ivl_15880 <= '0';
  tmp_ivl_15887 <= '0';
  tmp_ivl_15899 <= '0';
  tmp_ivl_15906 <= '0';
  tmp_ivl_15922 <= '0';
  tmp_ivl_15929 <= '0';
  tmp_ivl_15943 <= '0';
  tmp_ivl_15954 <= '0';
  tmp_ivl_15968 <= '0';
  tmp_ivl_15975 <= '0';
  tmp_ivl_15987 <= '0';
  tmp_ivl_15994 <= '0';
  tmp_ivl_16006 <= '0';
  tmp_ivl_16013 <= '0';
  tmp_ivl_16029 <= '0';
  tmp_ivl_16036 <= '0';
  tmp_ivl_1604 <= '0';
  tmp_ivl_16048 <= '0';
  tmp_ivl_16055 <= '0';
  tmp_ivl_16071 <= '0';
  tmp_ivl_16078 <= '0';
  tmp_ivl_16094 <= '0';
  tmp_ivl_16103 <= '0';
  tmp_ivl_16115 <= '0';
  tmp_ivl_16122 <= '0';
  tmp_ivl_16134 <= '0';
  tmp_ivl_16141 <= '0';
  tmp_ivl_1615 <= '0';
  tmp_ivl_16159 <= '0';
  tmp_ivl_16170 <= '0';
  tmp_ivl_16182 <= '0';
  tmp_ivl_16189 <= '0';
  tmp_ivl_16201 <= '0';
  tmp_ivl_16208 <= '0';
  tmp_ivl_16220 <= '0';
  tmp_ivl_16227 <= '0';
  tmp_ivl_16239 <= '0';
  tmp_ivl_16246 <= '0';
  tmp_ivl_16262 <= '0';
  tmp_ivl_16269 <= '0';
  tmp_ivl_16285 <= '0';
  tmp_ivl_16292 <= '0';
  tmp_ivl_16304 <= '0';
  tmp_ivl_16311 <= '0';
  tmp_ivl_16329 <= '0';
  tmp_ivl_1633 <= '0';
  tmp_ivl_16340 <= '0';
  tmp_ivl_16352 <= '0';
  tmp_ivl_16359 <= '0';
  tmp_ivl_16371 <= '0';
  tmp_ivl_16378 <= '0';
  tmp_ivl_16390 <= '0';
  tmp_ivl_16397 <= '0';
  tmp_ivl_16411 <= '0';
  tmp_ivl_16422 <= '0';
  tmp_ivl_16434 <= '0';
  tmp_ivl_1644 <= '0';
  tmp_ivl_16441 <= '0';
  tmp_ivl_16453 <= '0';
  tmp_ivl_16460 <= '0';
  tmp_ivl_16476 <= '0';
  tmp_ivl_16483 <= '0';
  tmp_ivl_16497 <= '0';
  tmp_ivl_165 <= '0';
  tmp_ivl_16508 <= '0';
  tmp_ivl_16524 <= '0';
  tmp_ivl_16531 <= '0';
  tmp_ivl_16543 <= '0';
  tmp_ivl_16550 <= '0';
  tmp_ivl_16562 <= '0';
  tmp_ivl_16569 <= '0';
  tmp_ivl_16587 <= '0';
  tmp_ivl_16598 <= '0';
  tmp_ivl_16610 <= '0';
  tmp_ivl_16617 <= '0';
  tmp_ivl_1662 <= '0';
  tmp_ivl_16629 <= '0';
  tmp_ivl_16636 <= '0';
  tmp_ivl_16648 <= '0';
  tmp_ivl_16655 <= '0';
  tmp_ivl_16667 <= '0';
  tmp_ivl_16674 <= '0';
  tmp_ivl_16686 <= '0';
  tmp_ivl_16693 <= '0';
  tmp_ivl_16711 <= '0';
  tmp_ivl_16722 <= '0';
  tmp_ivl_1673 <= '0';
  tmp_ivl_16738 <= '0';
  tmp_ivl_16745 <= '0';
  tmp_ivl_16757 <= '0';
  tmp_ivl_16764 <= '0';
  tmp_ivl_16776 <= '0';
  tmp_ivl_16783 <= '0';
  tmp_ivl_16797 <= '0';
  tmp_ivl_16808 <= '0';
  tmp_ivl_16824 <= '0';
  tmp_ivl_16831 <= '0';
  tmp_ivl_16843 <= '0';
  tmp_ivl_16850 <= '0';
  tmp_ivl_16862 <= '0';
  tmp_ivl_16869 <= '0';
  tmp_ivl_16885 <= '0';
  tmp_ivl_16892 <= '0';
  tmp_ivl_16904 <= '0';
  tmp_ivl_1691 <= '0';
  tmp_ivl_16911 <= '0';
  tmp_ivl_16927 <= '0';
  tmp_ivl_16934 <= '0';
  tmp_ivl_16950 <= '0';
  tmp_ivl_16959 <= '0';
  tmp_ivl_16975 <= '0';
  tmp_ivl_16982 <= '0';
  tmp_ivl_16994 <= '0';
  tmp_ivl_17001 <= '0';
  tmp_ivl_17017 <= '0';
  tmp_ivl_1702 <= '0';
  tmp_ivl_17024 <= '0';
  tmp_ivl_17036 <= '0';
  tmp_ivl_17043 <= '0';
  tmp_ivl_17059 <= '0';
  tmp_ivl_17066 <= '0';
  tmp_ivl_17078 <= '0';
  tmp_ivl_17085 <= '0';
  tmp_ivl_17101 <= '0';
  tmp_ivl_17108 <= '0';
  tmp_ivl_17122 <= '0';
  tmp_ivl_17133 <= '0';
  tmp_ivl_17147 <= '0';
  tmp_ivl_17158 <= '0';
  tmp_ivl_17174 <= '0';
  tmp_ivl_17181 <= '0';
  tmp_ivl_17193 <= '0';
  tmp_ivl_1720 <= '0';
  tmp_ivl_17200 <= '0';
  tmp_ivl_17212 <= '0';
  tmp_ivl_17219 <= '0';
  tmp_ivl_17235 <= '0';
  tmp_ivl_17242 <= '0';
  tmp_ivl_17256 <= '0';
  tmp_ivl_17267 <= '0';
  tmp_ivl_17281 <= '0';
  tmp_ivl_17288 <= '0';
  tmp_ivl_17300 <= '0';
  tmp_ivl_17307 <= '0';
  tmp_ivl_1731 <= '0';
  tmp_ivl_17319 <= '0';
  tmp_ivl_17326 <= '0';
  tmp_ivl_17342 <= '0';
  tmp_ivl_17349 <= '0';
  tmp_ivl_17361 <= '0';
  tmp_ivl_17368 <= '0';
  tmp_ivl_17386 <= '0';
  tmp_ivl_17397 <= '0';
  tmp_ivl_17409 <= '0';
  tmp_ivl_17416 <= '0';
  tmp_ivl_17428 <= '0';
  tmp_ivl_17435 <= '0';
  tmp_ivl_17447 <= '0';
  tmp_ivl_17454 <= '0';
  tmp_ivl_17466 <= '0';
  tmp_ivl_17473 <= '0';
  tmp_ivl_17489 <= '0';
  tmp_ivl_1749 <= '0';
  tmp_ivl_17496 <= '0';
  tmp_ivl_17510 <= '0';
  tmp_ivl_17521 <= '0';
  tmp_ivl_17537 <= '0';
  tmp_ivl_17544 <= '0';
  tmp_ivl_17556 <= '0';
  tmp_ivl_17563 <= '0';
  tmp_ivl_17575 <= '0';
  tmp_ivl_17582 <= '0';
  tmp_ivl_17598 <= '0';
  tmp_ivl_1760 <= '0';
  tmp_ivl_17605 <= '0';
  tmp_ivl_17621 <= '0';
  tmp_ivl_17630 <= '0';
  tmp_ivl_17642 <= '0';
  tmp_ivl_17649 <= '0';
  tmp_ivl_17661 <= '0';
  tmp_ivl_17668 <= '0';
  tmp_ivl_17684 <= '0';
  tmp_ivl_17691 <= '0';
  tmp_ivl_17703 <= '0';
  tmp_ivl_17710 <= '0';
  tmp_ivl_17726 <= '0';
  tmp_ivl_17733 <= '0';
  tmp_ivl_17749 <= '0';
  tmp_ivl_17756 <= '0';
  tmp_ivl_17768 <= '0';
  tmp_ivl_17775 <= '0';
  tmp_ivl_1778 <= '0';
  tmp_ivl_17791 <= '0';
  tmp_ivl_17798 <= '0';
  tmp_ivl_17812 <= '0';
  tmp_ivl_17823 <= '0';
  tmp_ivl_17837 <= '0';
  tmp_ivl_17848 <= '0';
  tmp_ivl_17864 <= '0';
  tmp_ivl_17871 <= '0';
  tmp_ivl_17883 <= '0';
  tmp_ivl_1789 <= '0';
  tmp_ivl_17890 <= '0';
  tmp_ivl_17902 <= '0';
  tmp_ivl_17909 <= '0';
  tmp_ivl_17925 <= '0';
  tmp_ivl_17932 <= '0';
  tmp_ivl_17946 <= '0';
  tmp_ivl_17953 <= '0';
  tmp_ivl_17965 <= '0';
  tmp_ivl_17972 <= '0';
  tmp_ivl_17984 <= '0';
  tmp_ivl_17991 <= '0';
  tmp_ivl_18009 <= '0';
  tmp_ivl_18020 <= '0';
  tmp_ivl_18032 <= '0';
  tmp_ivl_18039 <= '0';
  tmp_ivl_18051 <= '0';
  tmp_ivl_18058 <= '0';
  tmp_ivl_1807 <= '0';
  tmp_ivl_18070 <= '0';
  tmp_ivl_18077 <= '0';
  tmp_ivl_18089 <= '0';
  tmp_ivl_18096 <= '0';
  tmp_ivl_18112 <= '0';
  tmp_ivl_18119 <= '0';
  tmp_ivl_18133 <= '0';
  tmp_ivl_18144 <= '0';
  tmp_ivl_18160 <= '0';
  tmp_ivl_18167 <= '0';
  tmp_ivl_18179 <= '0';
  tmp_ivl_1818 <= '0';
  tmp_ivl_18186 <= '0';
  tmp_ivl_18198 <= '0';
  tmp_ivl_18205 <= '0';
  tmp_ivl_18221 <= '0';
  tmp_ivl_18228 <= '0';
  tmp_ivl_18244 <= '0';
  tmp_ivl_18253 <= '0';
  tmp_ivl_18269 <= '0';
  tmp_ivl_18276 <= '0';
  tmp_ivl_18288 <= '0';
  tmp_ivl_18295 <= '0';
  tmp_ivl_183 <= '0';
  tmp_ivl_18311 <= '0';
  tmp_ivl_18318 <= '0';
  tmp_ivl_18330 <= '0';
  tmp_ivl_18337 <= '0';
  tmp_ivl_18353 <= '0';
  tmp_ivl_1836 <= '0';
  tmp_ivl_18360 <= '0';
  tmp_ivl_18372 <= '0';
  tmp_ivl_18379 <= '0';
  tmp_ivl_18397 <= '0';
  tmp_ivl_18408 <= '0';
  tmp_ivl_18420 <= '0';
  tmp_ivl_18427 <= '0';
  tmp_ivl_18439 <= '0';
  tmp_ivl_18446 <= '0';
  tmp_ivl_18458 <= '0';
  tmp_ivl_18465 <= '0';
  tmp_ivl_1847 <= '0';
  tmp_ivl_18477 <= '0';
  tmp_ivl_18484 <= '0';
  tmp_ivl_18496 <= '0';
  tmp_ivl_18503 <= '0';
  tmp_ivl_18519 <= '0';
  tmp_ivl_18526 <= '0';
  tmp_ivl_18540 <= '0';
  tmp_ivl_18551 <= '0';
  tmp_ivl_18567 <= '0';
  tmp_ivl_18574 <= '0';
  tmp_ivl_18586 <= '0';
  tmp_ivl_18593 <= '0';
  tmp_ivl_18605 <= '0';
  tmp_ivl_18612 <= '0';
  tmp_ivl_18628 <= '0';
  tmp_ivl_18635 <= '0';
  tmp_ivl_18649 <= '0';
  tmp_ivl_1865 <= '0';
  tmp_ivl_18660 <= '0';
  tmp_ivl_18674 <= '0';
  tmp_ivl_18685 <= '0';
  tmp_ivl_18701 <= '0';
  tmp_ivl_18708 <= '0';
  tmp_ivl_18720 <= '0';
  tmp_ivl_18727 <= '0';
  tmp_ivl_18739 <= '0';
  tmp_ivl_18746 <= '0';
  tmp_ivl_1876 <= '0';
  tmp_ivl_18762 <= '0';
  tmp_ivl_18769 <= '0';
  tmp_ivl_18781 <= '0';
  tmp_ivl_18788 <= '0';
  tmp_ivl_18800 <= '0';
  tmp_ivl_18807 <= '0';
  tmp_ivl_18821 <= '0';
  tmp_ivl_18832 <= '0';
  tmp_ivl_18844 <= '0';
  tmp_ivl_18851 <= '0';
  tmp_ivl_18863 <= '0';
  tmp_ivl_18870 <= '0';
  tmp_ivl_18886 <= '0';
  tmp_ivl_18893 <= '0';
  tmp_ivl_18907 <= '0';
  tmp_ivl_18918 <= '0';
  tmp_ivl_18934 <= '0';
  tmp_ivl_1894 <= '0';
  tmp_ivl_18941 <= '0';
  tmp_ivl_18953 <= '0';
  tmp_ivl_18960 <= '0';
  tmp_ivl_18972 <= '0';
  tmp_ivl_18979 <= '0';
  tmp_ivl_18995 <= '0';
  tmp_ivl_19002 <= '0';
  tmp_ivl_19016 <= '0';
  tmp_ivl_19027 <= '0';
  tmp_ivl_19043 <= '0';
  tmp_ivl_1905 <= '0';
  tmp_ivl_19050 <= '0';
  tmp_ivl_19062 <= '0';
  tmp_ivl_19069 <= '0';
  tmp_ivl_19081 <= '0';
  tmp_ivl_19088 <= '0';
  tmp_ivl_19108 <= '0';
  tmp_ivl_19117 <= '0';
  tmp_ivl_19129 <= '0';
  tmp_ivl_19136 <= '0';
  tmp_ivl_19148 <= '0';
  tmp_ivl_19155 <= '0';
  tmp_ivl_19167 <= '0';
  tmp_ivl_19174 <= '0';
  tmp_ivl_19186 <= '0';
  tmp_ivl_19193 <= '0';
  tmp_ivl_19205 <= '0';
  tmp_ivl_19212 <= '0';
  tmp_ivl_19228 <= '0';
  tmp_ivl_1923 <= '0';
  tmp_ivl_19235 <= '0';
  tmp_ivl_19251 <= '0';
  tmp_ivl_19258 <= '0';
  tmp_ivl_19270 <= '0';
  tmp_ivl_19277 <= '0';
  tmp_ivl_19293 <= '0';
  tmp_ivl_19300 <= '0';
  tmp_ivl_19312 <= '0';
  tmp_ivl_19319 <= '0';
  tmp_ivl_19333 <= '0';
  tmp_ivl_1934 <= '0';
  tmp_ivl_19344 <= '0';
  tmp_ivl_19356 <= '0';
  tmp_ivl_19363 <= '0';
  tmp_ivl_19375 <= '0';
  tmp_ivl_19382 <= '0';
  tmp_ivl_19398 <= '0';
  tmp_ivl_194 <= '0';
  tmp_ivl_19405 <= '0';
  tmp_ivl_19419 <= '0';
  tmp_ivl_19426 <= '0';
  tmp_ivl_19438 <= '0';
  tmp_ivl_19445 <= '0';
  tmp_ivl_19457 <= '0';
  tmp_ivl_19464 <= '0';
  tmp_ivl_19480 <= '0';
  tmp_ivl_19487 <= '0';
  tmp_ivl_19499 <= '0';
  tmp_ivl_19506 <= '0';
  tmp_ivl_1952 <= '0';
  tmp_ivl_19520 <= '0';
  tmp_ivl_19531 <= '0';
  tmp_ivl_19543 <= '0';
  tmp_ivl_19550 <= '0';
  tmp_ivl_19562 <= '0';
  tmp_ivl_19569 <= '0';
  tmp_ivl_19585 <= '0';
  tmp_ivl_19592 <= '0';
  tmp_ivl_19606 <= '0';
  tmp_ivl_19617 <= '0';
  tmp_ivl_1963 <= '0';
  tmp_ivl_19633 <= '0';
  tmp_ivl_19640 <= '0';
  tmp_ivl_19652 <= '0';
  tmp_ivl_19659 <= '0';
  tmp_ivl_19671 <= '0';
  tmp_ivl_19678 <= '0';
  tmp_ivl_19694 <= '0';
  tmp_ivl_19701 <= '0';
  tmp_ivl_19717 <= '0';
  tmp_ivl_19726 <= '0';
  tmp_ivl_19738 <= '0';
  tmp_ivl_19745 <= '0';
  tmp_ivl_19757 <= '0';
  tmp_ivl_19764 <= '0';
  tmp_ivl_19780 <= '0';
  tmp_ivl_19787 <= '0';
  tmp_ivl_19803 <= '0';
  tmp_ivl_1981 <= '0';
  tmp_ivl_19810 <= '0';
  tmp_ivl_19822 <= '0';
  tmp_ivl_19829 <= '0';
  tmp_ivl_19845 <= '0';
  tmp_ivl_19852 <= '0';
  tmp_ivl_19864 <= '0';
  tmp_ivl_19871 <= '0';
  tmp_ivl_19887 <= '0';
  tmp_ivl_19894 <= '0';
  tmp_ivl_19906 <= '0';
  tmp_ivl_19913 <= '0';
  tmp_ivl_1992 <= '0';
  tmp_ivl_19929 <= '0';
  tmp_ivl_19936 <= '0';
  tmp_ivl_19950 <= '0';
  tmp_ivl_19961 <= '0';
  tmp_ivl_19973 <= '0';
  tmp_ivl_19980 <= '0';
  tmp_ivl_19992 <= '0';
  tmp_ivl_19999 <= '0';
  tmp_ivl_20 <= '0';
  tmp_ivl_20015 <= '0';
  tmp_ivl_20022 <= '0';
  tmp_ivl_20034 <= '0';
  tmp_ivl_20041 <= '0';
  tmp_ivl_20057 <= '0';
  tmp_ivl_20064 <= '0';
  tmp_ivl_20078 <= '0';
  tmp_ivl_20089 <= '0';
  tmp_ivl_2010 <= '0';
  tmp_ivl_20105 <= '0';
  tmp_ivl_20112 <= '0';
  tmp_ivl_20124 <= '0';
  tmp_ivl_20131 <= '0';
  tmp_ivl_20143 <= '0';
  tmp_ivl_20150 <= '0';
  tmp_ivl_20166 <= '0';
  tmp_ivl_20173 <= '0';
  tmp_ivl_20185 <= '0';
  tmp_ivl_20192 <= '0';
  tmp_ivl_20208 <= '0';
  tmp_ivl_2021 <= '0';
  tmp_ivl_20215 <= '0';
  tmp_ivl_20229 <= '0';
  tmp_ivl_20240 <= '0';
  tmp_ivl_20252 <= '0';
  tmp_ivl_20259 <= '0';
  tmp_ivl_20271 <= '0';
  tmp_ivl_20278 <= '0';
  tmp_ivl_20294 <= '0';
  tmp_ivl_20301 <= '0';
  tmp_ivl_20315 <= '0';
  tmp_ivl_20326 <= '0';
  tmp_ivl_20342 <= '0';
  tmp_ivl_20349 <= '0';
  tmp_ivl_20361 <= '0';
  tmp_ivl_20368 <= '0';
  tmp_ivl_20380 <= '0';
  tmp_ivl_20387 <= '0';
  tmp_ivl_2039 <= '0';
  tmp_ivl_20403 <= '0';
  tmp_ivl_20410 <= '0';
  tmp_ivl_20426 <= '0';
  tmp_ivl_20435 <= '0';
  tmp_ivl_20447 <= '0';
  tmp_ivl_20454 <= '0';
  tmp_ivl_20466 <= '0';
  tmp_ivl_20473 <= '0';
  tmp_ivl_20489 <= '0';
  tmp_ivl_20496 <= '0';
  tmp_ivl_2050 <= '0';
  tmp_ivl_20508 <= '0';
  tmp_ivl_20515 <= '0';
  tmp_ivl_20531 <= '0';
  tmp_ivl_20538 <= '0';
  tmp_ivl_20554 <= '0';
  tmp_ivl_20561 <= '0';
  tmp_ivl_20573 <= '0';
  tmp_ivl_20580 <= '0';
  tmp_ivl_20596 <= '0';
  tmp_ivl_20603 <= '0';
  tmp_ivl_20615 <= '0';
  tmp_ivl_20622 <= '0';
  tmp_ivl_20638 <= '0';
  tmp_ivl_20645 <= '0';
  tmp_ivl_20657 <= '0';
  tmp_ivl_20664 <= '0';
  tmp_ivl_2068 <= '0';
  tmp_ivl_20680 <= '0';
  tmp_ivl_20687 <= '0';
  tmp_ivl_20701 <= '0';
  tmp_ivl_20712 <= '0';
  tmp_ivl_20724 <= '0';
  tmp_ivl_20731 <= '0';
  tmp_ivl_20743 <= '0';
  tmp_ivl_20750 <= '0';
  tmp_ivl_20766 <= '0';
  tmp_ivl_20773 <= '0';
  tmp_ivl_20785 <= '0';
  tmp_ivl_2079 <= '0';
  tmp_ivl_20792 <= '0';
  tmp_ivl_20808 <= '0';
  tmp_ivl_20815 <= '0';
  tmp_ivl_20829 <= '0';
  tmp_ivl_20840 <= '0';
  tmp_ivl_20856 <= '0';
  tmp_ivl_20863 <= '0';
  tmp_ivl_20875 <= '0';
  tmp_ivl_20882 <= '0';
  tmp_ivl_20894 <= '0';
  tmp_ivl_20901 <= '0';
  tmp_ivl_20917 <= '0';
  tmp_ivl_20924 <= '0';
  tmp_ivl_20936 <= '0';
  tmp_ivl_20943 <= '0';
  tmp_ivl_20959 <= '0';
  tmp_ivl_20966 <= '0';
  tmp_ivl_2097 <= '0';
  tmp_ivl_20982 <= '0';
  tmp_ivl_20991 <= '0';
  tmp_ivl_21003 <= '0';
  tmp_ivl_21010 <= '0';
  tmp_ivl_21022 <= '0';
  tmp_ivl_21029 <= '0';
  tmp_ivl_21041 <= '0';
  tmp_ivl_21048 <= '0';
  tmp_ivl_21060 <= '0';
  tmp_ivl_21067 <= '0';
  tmp_ivl_2108 <= '0';
  tmp_ivl_21083 <= '0';
  tmp_ivl_21090 <= '0';
  tmp_ivl_21106 <= '0';
  tmp_ivl_21113 <= '0';
  tmp_ivl_21125 <= '0';
  tmp_ivl_21132 <= '0';
  tmp_ivl_21148 <= '0';
  tmp_ivl_21155 <= '0';
  tmp_ivl_21167 <= '0';
  tmp_ivl_21174 <= '0';
  tmp_ivl_21190 <= '0';
  tmp_ivl_21197 <= '0';
  tmp_ivl_212 <= '0';
  tmp_ivl_21211 <= '0';
  tmp_ivl_21222 <= '0';
  tmp_ivl_21234 <= '0';
  tmp_ivl_21241 <= '0';
  tmp_ivl_21253 <= '0';
  tmp_ivl_2126 <= '0';
  tmp_ivl_21260 <= '0';
  tmp_ivl_21276 <= '0';
  tmp_ivl_21283 <= '0';
  tmp_ivl_21295 <= '0';
  tmp_ivl_21302 <= '0';
  tmp_ivl_21318 <= '0';
  tmp_ivl_21325 <= '0';
  tmp_ivl_21337 <= '0';
  tmp_ivl_21344 <= '0';
  tmp_ivl_21360 <= '0';
  tmp_ivl_21367 <= '0';
  tmp_ivl_2137 <= '0';
  tmp_ivl_21381 <= '0';
  tmp_ivl_21388 <= '0';
  tmp_ivl_21400 <= '0';
  tmp_ivl_21407 <= '0';
  tmp_ivl_21419 <= '0';
  tmp_ivl_21426 <= '0';
  tmp_ivl_21442 <= '0';
  tmp_ivl_21449 <= '0';
  tmp_ivl_21461 <= '0';
  tmp_ivl_21468 <= '0';
  tmp_ivl_21484 <= '0';
  tmp_ivl_21491 <= '0';
  tmp_ivl_21505 <= '0';
  tmp_ivl_21516 <= '0';
  tmp_ivl_21528 <= '0';
  tmp_ivl_21535 <= '0';
  tmp_ivl_21547 <= '0';
  tmp_ivl_2155 <= '0';
  tmp_ivl_21554 <= '0';
  tmp_ivl_21570 <= '0';
  tmp_ivl_21577 <= '0';
  tmp_ivl_21589 <= '0';
  tmp_ivl_21596 <= '0';
  tmp_ivl_21612 <= '0';
  tmp_ivl_21619 <= '0';
  tmp_ivl_21631 <= '0';
  tmp_ivl_21638 <= '0';
  tmp_ivl_21654 <= '0';
  tmp_ivl_2166 <= '0';
  tmp_ivl_21661 <= '0';
  tmp_ivl_21675 <= '0';
  tmp_ivl_21686 <= '0';
  tmp_ivl_21702 <= '0';
  tmp_ivl_21709 <= '0';
  tmp_ivl_21721 <= '0';
  tmp_ivl_21728 <= '0';
  tmp_ivl_21740 <= '0';
  tmp_ivl_21747 <= '0';
  tmp_ivl_21763 <= '0';
  tmp_ivl_21770 <= '0';
  tmp_ivl_21782 <= '0';
  tmp_ivl_21789 <= '0';
  tmp_ivl_21805 <= '0';
  tmp_ivl_21812 <= '0';
  tmp_ivl_21828 <= '0';
  tmp_ivl_21837 <= '0';
  tmp_ivl_2184 <= '0';
  tmp_ivl_21849 <= '0';
  tmp_ivl_21856 <= '0';
  tmp_ivl_21868 <= '0';
  tmp_ivl_21875 <= '0';
  tmp_ivl_21891 <= '0';
  tmp_ivl_21898 <= '0';
  tmp_ivl_21910 <= '0';
  tmp_ivl_21917 <= '0';
  tmp_ivl_21933 <= '0';
  tmp_ivl_21940 <= '0';
  tmp_ivl_2195 <= '0';
  tmp_ivl_21956 <= '0';
  tmp_ivl_21963 <= '0';
  tmp_ivl_21975 <= '0';
  tmp_ivl_21982 <= '0';
  tmp_ivl_21998 <= '0';
  tmp_ivl_22005 <= '0';
  tmp_ivl_22017 <= '0';
  tmp_ivl_22024 <= '0';
  tmp_ivl_22040 <= '0';
  tmp_ivl_22047 <= '0';
  tmp_ivl_22059 <= '0';
  tmp_ivl_22066 <= '0';
  tmp_ivl_22082 <= '0';
  tmp_ivl_22089 <= '0';
  tmp_ivl_22103 <= '0';
  tmp_ivl_22114 <= '0';
  tmp_ivl_22126 <= '0';
  tmp_ivl_2213 <= '0';
  tmp_ivl_22133 <= '0';
  tmp_ivl_22145 <= '0';
  tmp_ivl_22152 <= '0';
  tmp_ivl_22168 <= '0';
  tmp_ivl_22175 <= '0';
  tmp_ivl_22187 <= '0';
  tmp_ivl_22194 <= '0';
  tmp_ivl_22210 <= '0';
  tmp_ivl_22217 <= '0';
  tmp_ivl_22229 <= '0';
  tmp_ivl_22236 <= '0';
  tmp_ivl_2224 <= '0';
  tmp_ivl_22252 <= '0';
  tmp_ivl_22259 <= '0';
  tmp_ivl_22273 <= '0';
  tmp_ivl_22284 <= '0';
  tmp_ivl_223 <= '0';
  tmp_ivl_22300 <= '0';
  tmp_ivl_22307 <= '0';
  tmp_ivl_22319 <= '0';
  tmp_ivl_22326 <= '0';
  tmp_ivl_22338 <= '0';
  tmp_ivl_22345 <= '0';
  tmp_ivl_22361 <= '0';
  tmp_ivl_22368 <= '0';
  tmp_ivl_22380 <= '0';
  tmp_ivl_22387 <= '0';
  tmp_ivl_22403 <= '0';
  tmp_ivl_22410 <= '0';
  tmp_ivl_2242 <= '0';
  tmp_ivl_22422 <= '0';
  tmp_ivl_22429 <= '0';
  tmp_ivl_22445 <= '0';
  tmp_ivl_22452 <= '0';
  tmp_ivl_22466 <= '0';
  tmp_ivl_22477 <= '0';
  tmp_ivl_22489 <= '0';
  tmp_ivl_22496 <= '0';
  tmp_ivl_22508 <= '0';
  tmp_ivl_22515 <= '0';
  tmp_ivl_2253 <= '0';
  tmp_ivl_22531 <= '0';
  tmp_ivl_22538 <= '0';
  tmp_ivl_22550 <= '0';
  tmp_ivl_22557 <= '0';
  tmp_ivl_22573 <= '0';
  tmp_ivl_22580 <= '0';
  tmp_ivl_22594 <= '0';
  tmp_ivl_22605 <= '0';
  tmp_ivl_22621 <= '0';
  tmp_ivl_22628 <= '0';
  tmp_ivl_22640 <= '0';
  tmp_ivl_22647 <= '0';
  tmp_ivl_22659 <= '0';
  tmp_ivl_22666 <= '0';
  tmp_ivl_22682 <= '0';
  tmp_ivl_22689 <= '0';
  tmp_ivl_22701 <= '0';
  tmp_ivl_22708 <= '0';
  tmp_ivl_2271 <= '0';
  tmp_ivl_22724 <= '0';
  tmp_ivl_22731 <= '0';
  tmp_ivl_22743 <= '0';
  tmp_ivl_22750 <= '0';
  tmp_ivl_22766 <= '0';
  tmp_ivl_22775 <= '0';
  tmp_ivl_22787 <= '0';
  tmp_ivl_22794 <= '0';
  tmp_ivl_22806 <= '0';
  tmp_ivl_22813 <= '0';
  tmp_ivl_2282 <= '0';
  tmp_ivl_22829 <= '0';
  tmp_ivl_22836 <= '0';
  tmp_ivl_22848 <= '0';
  tmp_ivl_22855 <= '0';
  tmp_ivl_22871 <= '0';
  tmp_ivl_22878 <= '0';
  tmp_ivl_22894 <= '0';
  tmp_ivl_22901 <= '0';
  tmp_ivl_22913 <= '0';
  tmp_ivl_22920 <= '0';
  tmp_ivl_22936 <= '0';
  tmp_ivl_22943 <= '0';
  tmp_ivl_22955 <= '0';
  tmp_ivl_22962 <= '0';
  tmp_ivl_22978 <= '0';
  tmp_ivl_22985 <= '0';
  tmp_ivl_22999 <= '0';
  tmp_ivl_2300 <= '0';
  tmp_ivl_23010 <= '0';
  tmp_ivl_23022 <= '0';
  tmp_ivl_23029 <= '0';
  tmp_ivl_23041 <= '0';
  tmp_ivl_23048 <= '0';
  tmp_ivl_23064 <= '0';
  tmp_ivl_23071 <= '0';
  tmp_ivl_23083 <= '0';
  tmp_ivl_23090 <= '0';
  tmp_ivl_23106 <= '0';
  tmp_ivl_2311 <= '0';
  tmp_ivl_23113 <= '0';
  tmp_ivl_23125 <= '0';
  tmp_ivl_23132 <= '0';
  tmp_ivl_23148 <= '0';
  tmp_ivl_23155 <= '0';
  tmp_ivl_23169 <= '0';
  tmp_ivl_23176 <= '0';
  tmp_ivl_23188 <= '0';
  tmp_ivl_23195 <= '0';
  tmp_ivl_23207 <= '0';
  tmp_ivl_23214 <= '0';
  tmp_ivl_23230 <= '0';
  tmp_ivl_23237 <= '0';
  tmp_ivl_23249 <= '0';
  tmp_ivl_23256 <= '0';
  tmp_ivl_23272 <= '0';
  tmp_ivl_23279 <= '0';
  tmp_ivl_2329 <= '0';
  tmp_ivl_23293 <= '0';
  tmp_ivl_23304 <= '0';
  tmp_ivl_23316 <= '0';
  tmp_ivl_23323 <= '0';
  tmp_ivl_23335 <= '0';
  tmp_ivl_23342 <= '0';
  tmp_ivl_23358 <= '0';
  tmp_ivl_23365 <= '0';
  tmp_ivl_23377 <= '0';
  tmp_ivl_23384 <= '0';
  tmp_ivl_2340 <= '0';
  tmp_ivl_23400 <= '0';
  tmp_ivl_23407 <= '0';
  tmp_ivl_23419 <= '0';
  tmp_ivl_23426 <= '0';
  tmp_ivl_23442 <= '0';
  tmp_ivl_23449 <= '0';
  tmp_ivl_23463 <= '0';
  tmp_ivl_23474 <= '0';
  tmp_ivl_23490 <= '0';
  tmp_ivl_23497 <= '0';
  tmp_ivl_23509 <= '0';
  tmp_ivl_23516 <= '0';
  tmp_ivl_23528 <= '0';
  tmp_ivl_23535 <= '0';
  tmp_ivl_23551 <= '0';
  tmp_ivl_23558 <= '0';
  tmp_ivl_23570 <= '0';
  tmp_ivl_23577 <= '0';
  tmp_ivl_2358 <= '0';
  tmp_ivl_23593 <= '0';
  tmp_ivl_23600 <= '0';
  tmp_ivl_23612 <= '0';
  tmp_ivl_23619 <= '0';
  tmp_ivl_23635 <= '0';
  tmp_ivl_23642 <= '0';
  tmp_ivl_23658 <= '0';
  tmp_ivl_23667 <= '0';
  tmp_ivl_23679 <= '0';
  tmp_ivl_23686 <= '0';
  tmp_ivl_2369 <= '0';
  tmp_ivl_23698 <= '0';
  tmp_ivl_23705 <= '0';
  tmp_ivl_23721 <= '0';
  tmp_ivl_23728 <= '0';
  tmp_ivl_23740 <= '0';
  tmp_ivl_23747 <= '0';
  tmp_ivl_23763 <= '0';
  tmp_ivl_23770 <= '0';
  tmp_ivl_23782 <= '0';
  tmp_ivl_23789 <= '0';
  tmp_ivl_23805 <= '0';
  tmp_ivl_23812 <= '0';
  tmp_ivl_23828 <= '0';
  tmp_ivl_23835 <= '0';
  tmp_ivl_23847 <= '0';
  tmp_ivl_23854 <= '0';
  tmp_ivl_2387 <= '0';
  tmp_ivl_23870 <= '0';
  tmp_ivl_23877 <= '0';
  tmp_ivl_23889 <= '0';
  tmp_ivl_23896 <= '0';
  tmp_ivl_23912 <= '0';
  tmp_ivl_23919 <= '0';
  tmp_ivl_23931 <= '0';
  tmp_ivl_23938 <= '0';
  tmp_ivl_23954 <= '0';
  tmp_ivl_23961 <= '0';
  tmp_ivl_23975 <= '0';
  tmp_ivl_2398 <= '0';
  tmp_ivl_23986 <= '0';
  tmp_ivl_23998 <= '0';
  tmp_ivl_24005 <= '0';
  tmp_ivl_24017 <= '0';
  tmp_ivl_24024 <= '0';
  tmp_ivl_24040 <= '0';
  tmp_ivl_24047 <= '0';
  tmp_ivl_24059 <= '0';
  tmp_ivl_24066 <= '0';
  tmp_ivl_24082 <= '0';
  tmp_ivl_24089 <= '0';
  tmp_ivl_241 <= '0';
  tmp_ivl_24103 <= '0';
  tmp_ivl_24114 <= '0';
  tmp_ivl_24130 <= '0';
  tmp_ivl_24137 <= '0';
  tmp_ivl_24149 <= '0';
  tmp_ivl_24156 <= '0';
  tmp_ivl_2416 <= '0';
  tmp_ivl_24168 <= '0';
  tmp_ivl_24175 <= '0';
  tmp_ivl_24191 <= '0';
  tmp_ivl_24198 <= '0';
  tmp_ivl_24210 <= '0';
  tmp_ivl_24217 <= '0';
  tmp_ivl_24233 <= '0';
  tmp_ivl_24240 <= '0';
  tmp_ivl_24256 <= '0';
  tmp_ivl_24265 <= '0';
  tmp_ivl_2427 <= '0';
  tmp_ivl_24277 <= '0';
  tmp_ivl_24284 <= '0';
  tmp_ivl_24296 <= '0';
  tmp_ivl_24303 <= '0';
  tmp_ivl_24319 <= '0';
  tmp_ivl_24326 <= '0';
  tmp_ivl_24338 <= '0';
  tmp_ivl_24345 <= '0';
  tmp_ivl_24361 <= '0';
  tmp_ivl_24368 <= '0';
  tmp_ivl_24380 <= '0';
  tmp_ivl_24387 <= '0';
  tmp_ivl_24403 <= '0';
  tmp_ivl_24410 <= '0';
  tmp_ivl_24426 <= '0';
  tmp_ivl_24433 <= '0';
  tmp_ivl_24445 <= '0';
  tmp_ivl_2445 <= '0';
  tmp_ivl_24452 <= '0';
  tmp_ivl_24468 <= '0';
  tmp_ivl_24475 <= '0';
  tmp_ivl_24487 <= '0';
  tmp_ivl_24494 <= '0';
  tmp_ivl_24510 <= '0';
  tmp_ivl_24517 <= '0';
  tmp_ivl_24531 <= '0';
  tmp_ivl_24542 <= '0';
  tmp_ivl_24554 <= '0';
  tmp_ivl_2456 <= '0';
  tmp_ivl_24561 <= '0';
  tmp_ivl_24573 <= '0';
  tmp_ivl_24580 <= '0';
  tmp_ivl_24596 <= '0';
  tmp_ivl_24603 <= '0';
  tmp_ivl_24615 <= '0';
  tmp_ivl_24622 <= '0';
  tmp_ivl_24638 <= '0';
  tmp_ivl_24645 <= '0';
  tmp_ivl_24659 <= '0';
  tmp_ivl_24670 <= '0';
  tmp_ivl_24686 <= '0';
  tmp_ivl_24693 <= '0';
  tmp_ivl_24705 <= '0';
  tmp_ivl_24712 <= '0';
  tmp_ivl_24724 <= '0';
  tmp_ivl_24731 <= '0';
  tmp_ivl_2474 <= '0';
  tmp_ivl_24747 <= '0';
  tmp_ivl_24754 <= '0';
  tmp_ivl_24766 <= '0';
  tmp_ivl_24773 <= '0';
  tmp_ivl_24789 <= '0';
  tmp_ivl_24796 <= '0';
  tmp_ivl_24810 <= '0';
  tmp_ivl_24821 <= '0';
  tmp_ivl_24833 <= '0';
  tmp_ivl_24840 <= '0';
  tmp_ivl_2485 <= '0';
  tmp_ivl_24852 <= '0';
  tmp_ivl_24859 <= '0';
  tmp_ivl_24875 <= '0';
  tmp_ivl_24882 <= '0';
  tmp_ivl_24894 <= '0';
  tmp_ivl_24901 <= '0';
  tmp_ivl_24917 <= '0';
  tmp_ivl_24924 <= '0';
  tmp_ivl_24936 <= '0';
  tmp_ivl_24943 <= '0';
  tmp_ivl_24959 <= '0';
  tmp_ivl_24966 <= '0';
  tmp_ivl_24980 <= '0';
  tmp_ivl_24991 <= '0';
  tmp_ivl_25007 <= '0';
  tmp_ivl_25014 <= '0';
  tmp_ivl_25026 <= '0';
  tmp_ivl_2503 <= '0';
  tmp_ivl_25033 <= '0';
  tmp_ivl_25045 <= '0';
  tmp_ivl_25052 <= '0';
  tmp_ivl_25068 <= '0';
  tmp_ivl_25075 <= '0';
  tmp_ivl_25087 <= '0';
  tmp_ivl_25094 <= '0';
  tmp_ivl_25110 <= '0';
  tmp_ivl_25117 <= '0';
  tmp_ivl_25129 <= '0';
  tmp_ivl_25136 <= '0';
  tmp_ivl_2514 <= '0';
  tmp_ivl_25152 <= '0';
  tmp_ivl_25159 <= '0';
  tmp_ivl_25175 <= '0';
  tmp_ivl_25184 <= '0';
  tmp_ivl_25196 <= '0';
  tmp_ivl_252 <= '0';
  tmp_ivl_25203 <= '0';
  tmp_ivl_25215 <= '0';
  tmp_ivl_25222 <= '0';
  tmp_ivl_25238 <= '0';
  tmp_ivl_25245 <= '0';
  tmp_ivl_25257 <= '0';
  tmp_ivl_25264 <= '0';
  tmp_ivl_25280 <= '0';
  tmp_ivl_25287 <= '0';
  tmp_ivl_25299 <= '0';
  tmp_ivl_25306 <= '0';
  tmp_ivl_2532 <= '0';
  tmp_ivl_25322 <= '0';
  tmp_ivl_25329 <= '0';
  tmp_ivl_25345 <= '0';
  tmp_ivl_25352 <= '0';
  tmp_ivl_25364 <= '0';
  tmp_ivl_25371 <= '0';
  tmp_ivl_25387 <= '0';
  tmp_ivl_25394 <= '0';
  tmp_ivl_25406 <= '0';
  tmp_ivl_25413 <= '0';
  tmp_ivl_25429 <= '0';
  tmp_ivl_2543 <= '0';
  tmp_ivl_25436 <= '0';
  tmp_ivl_25448 <= '0';
  tmp_ivl_25455 <= '0';
  tmp_ivl_25471 <= '0';
  tmp_ivl_25480 <= '0';
  tmp_ivl_25494 <= '0';
  tmp_ivl_25505 <= '0';
  tmp_ivl_25517 <= '0';
  tmp_ivl_25524 <= '0';
  tmp_ivl_25536 <= '0';
  tmp_ivl_25545 <= '0';
  tmp_ivl_25559 <= '0';
  tmp_ivl_25570 <= '0';
  tmp_ivl_25582 <= '0';
  tmp_ivl_25589 <= '0';
  tmp_ivl_25601 <= '0';
  tmp_ivl_25608 <= '0';
  tmp_ivl_2561 <= '0';
  tmp_ivl_25620 <= '0';
  tmp_ivl_25629 <= '0';
  tmp_ivl_25643 <= '0';
  tmp_ivl_25654 <= '0';
  tmp_ivl_25666 <= '0';
  tmp_ivl_25673 <= '0';
  tmp_ivl_25685 <= '0';
  tmp_ivl_25692 <= '0';
  tmp_ivl_25708 <= '0';
  tmp_ivl_25717 <= '0';
  tmp_ivl_2572 <= '0';
  tmp_ivl_25731 <= '0';
  tmp_ivl_25742 <= '0';
  tmp_ivl_25754 <= '0';
  tmp_ivl_25761 <= '0';
  tmp_ivl_25773 <= '0';
  tmp_ivl_25782 <= '0';
  tmp_ivl_25796 <= '0';
  tmp_ivl_25807 <= '0';
  tmp_ivl_25819 <= '0';
  tmp_ivl_25826 <= '0';
  tmp_ivl_25838 <= '0';
  tmp_ivl_25845 <= '0';
  tmp_ivl_25857 <= '0';
  tmp_ivl_25866 <= '0';
  tmp_ivl_25880 <= '0';
  tmp_ivl_25891 <= '0';
  tmp_ivl_2590 <= '0';
  tmp_ivl_25903 <= '0';
  tmp_ivl_25910 <= '0';
  tmp_ivl_25922 <= '0';
  tmp_ivl_25929 <= '0';
  tmp_ivl_25945 <= '0';
  tmp_ivl_25954 <= '0';
  tmp_ivl_25968 <= '0';
  tmp_ivl_25979 <= '0';
  tmp_ivl_25991 <= '0';
  tmp_ivl_25998 <= '0';
  tmp_ivl_2601 <= '0';
  tmp_ivl_26010 <= '0';
  tmp_ivl_26019 <= '0';
  tmp_ivl_26033 <= '0';
  tmp_ivl_26044 <= '0';
  tmp_ivl_26056 <= '0';
  tmp_ivl_26063 <= '0';
  tmp_ivl_26075 <= '0';
  tmp_ivl_26084 <= '0';
  tmp_ivl_26098 <= '0';
  tmp_ivl_26109 <= '0';
  tmp_ivl_26121 <= '0';
  tmp_ivl_26128 <= '0';
  tmp_ivl_26140 <= '0';
  tmp_ivl_26147 <= '0';
  tmp_ivl_26159 <= '0';
  tmp_ivl_26166 <= '0';
  tmp_ivl_26182 <= '0';
  tmp_ivl_2619 <= '0';
  tmp_ivl_26191 <= '0';
  tmp_ivl_26205 <= '0';
  tmp_ivl_26216 <= '0';
  tmp_ivl_26228 <= '0';
  tmp_ivl_26235 <= '0';
  tmp_ivl_26247 <= '0';
  tmp_ivl_26256 <= '0';
  tmp_ivl_26270 <= '0';
  tmp_ivl_26281 <= '0';
  tmp_ivl_26293 <= '0';
  tmp_ivl_2630 <= '0';
  tmp_ivl_26300 <= '0';
  tmp_ivl_26312 <= '0';
  tmp_ivl_26321 <= '0';
  tmp_ivl_26335 <= '0';
  tmp_ivl_26346 <= '0';
  tmp_ivl_26358 <= '0';
  tmp_ivl_26365 <= '0';
  tmp_ivl_26377 <= '0';
  tmp_ivl_26384 <= '0';
  tmp_ivl_26396 <= '0';
  tmp_ivl_26403 <= '0';
  tmp_ivl_26419 <= '0';
  tmp_ivl_26428 <= '0';
  tmp_ivl_26442 <= '0';
  tmp_ivl_26453 <= '0';
  tmp_ivl_26465 <= '0';
  tmp_ivl_26472 <= '0';
  tmp_ivl_2648 <= '0';
  tmp_ivl_26484 <= '0';
  tmp_ivl_26493 <= '0';
  tmp_ivl_26507 <= '0';
  tmp_ivl_26518 <= '0';
  tmp_ivl_26530 <= '0';
  tmp_ivl_26537 <= '0';
  tmp_ivl_26549 <= '0';
  tmp_ivl_26556 <= '0';
  tmp_ivl_26568 <= '0';
  tmp_ivl_26577 <= '0';
  tmp_ivl_2659 <= '0';
  tmp_ivl_26591 <= '0';
  tmp_ivl_26602 <= '0';
  tmp_ivl_26614 <= '0';
  tmp_ivl_26621 <= '0';
  tmp_ivl_26633 <= '0';
  tmp_ivl_26640 <= '0';
  tmp_ivl_26656 <= '0';
  tmp_ivl_26665 <= '0';
  tmp_ivl_26679 <= '0';
  tmp_ivl_26690 <= '0';
  tmp_ivl_26702 <= '0';
  tmp_ivl_26709 <= '0';
  tmp_ivl_26721 <= '0';
  tmp_ivl_26730 <= '0';
  tmp_ivl_26744 <= '0';
  tmp_ivl_26755 <= '0';
  tmp_ivl_26767 <= '0';
  tmp_ivl_2677 <= '0';
  tmp_ivl_26774 <= '0';
  tmp_ivl_26786 <= '0';
  tmp_ivl_26793 <= '0';
  tmp_ivl_26805 <= '0';
  tmp_ivl_26814 <= '0';
  tmp_ivl_26828 <= '0';
  tmp_ivl_26839 <= '0';
  tmp_ivl_26851 <= '0';
  tmp_ivl_26858 <= '0';
  tmp_ivl_26870 <= '0';
  tmp_ivl_26877 <= '0';
  tmp_ivl_2688 <= '0';
  tmp_ivl_26893 <= '0';
  tmp_ivl_26902 <= '0';
  tmp_ivl_26916 <= '0';
  tmp_ivl_26927 <= '0';
  tmp_ivl_26939 <= '0';
  tmp_ivl_26946 <= '0';
  tmp_ivl_26958 <= '0';
  tmp_ivl_26967 <= '0';
  tmp_ivl_26981 <= '0';
  tmp_ivl_26992 <= '0';
  tmp_ivl_270 <= '0';
  tmp_ivl_27004 <= '0';
  tmp_ivl_27011 <= '0';
  tmp_ivl_27023 <= '0';
  tmp_ivl_27032 <= '0';
  tmp_ivl_27046 <= '0';
  tmp_ivl_27057 <= '0';
  tmp_ivl_2706 <= '0';
  tmp_ivl_27069 <= '0';
  tmp_ivl_27076 <= '0';
  tmp_ivl_27088 <= '0';
  tmp_ivl_27095 <= '0';
  tmp_ivl_27107 <= '0';
  tmp_ivl_27114 <= '0';
  tmp_ivl_27130 <= '0';
  tmp_ivl_27139 <= '0';
  tmp_ivl_27153 <= '0';
  tmp_ivl_27164 <= '0';
  tmp_ivl_2717 <= '0';
  tmp_ivl_27176 <= '0';
  tmp_ivl_27183 <= '0';
  tmp_ivl_27195 <= '0';
  tmp_ivl_27202 <= '0';
  tmp_ivl_27214 <= '0';
  tmp_ivl_27223 <= '0';
  tmp_ivl_27237 <= '0';
  tmp_ivl_27248 <= '0';
  tmp_ivl_27260 <= '0';
  tmp_ivl_27267 <= '0';
  tmp_ivl_27279 <= '0';
  tmp_ivl_27286 <= '0';
  tmp_ivl_27302 <= '0';
  tmp_ivl_27311 <= '0';
  tmp_ivl_27325 <= '0';
  tmp_ivl_27336 <= '0';
  tmp_ivl_27348 <= '0';
  tmp_ivl_2735 <= '0';
  tmp_ivl_27355 <= '0';
  tmp_ivl_27367 <= '0';
  tmp_ivl_27374 <= '0';
  tmp_ivl_27386 <= '0';
  tmp_ivl_27395 <= '0';
  tmp_ivl_27409 <= '0';
  tmp_ivl_27420 <= '0';
  tmp_ivl_27432 <= '0';
  tmp_ivl_27439 <= '0';
  tmp_ivl_27451 <= '0';
  tmp_ivl_27458 <= '0';
  tmp_ivl_2746 <= '0';
  tmp_ivl_27474 <= '0';
  tmp_ivl_27483 <= '0';
  tmp_ivl_27497 <= '0';
  tmp_ivl_27508 <= '0';
  tmp_ivl_27520 <= '0';
  tmp_ivl_27527 <= '0';
  tmp_ivl_27539 <= '0';
  tmp_ivl_27548 <= '0';
  tmp_ivl_27562 <= '0';
  tmp_ivl_27573 <= '0';
  tmp_ivl_27585 <= '0';
  tmp_ivl_27592 <= '0';
  tmp_ivl_27604 <= '0';
  tmp_ivl_27611 <= '0';
  tmp_ivl_27623 <= '0';
  tmp_ivl_27630 <= '0';
  tmp_ivl_2764 <= '0';
  tmp_ivl_27646 <= '0';
  tmp_ivl_27653 <= '0';
  tmp_ivl_27665 <= '0';
  tmp_ivl_27674 <= '0';
  tmp_ivl_27688 <= '0';
  tmp_ivl_27699 <= '0';
  tmp_ivl_27711 <= '0';
  tmp_ivl_27718 <= '0';
  tmp_ivl_27730 <= '0';
  tmp_ivl_27737 <= '0';
  tmp_ivl_2775 <= '0';
  tmp_ivl_27753 <= '0';
  tmp_ivl_27760 <= '0';
  tmp_ivl_27772 <= '0';
  tmp_ivl_27781 <= '0';
  tmp_ivl_27795 <= '0';
  tmp_ivl_27806 <= '0';
  tmp_ivl_27818 <= '0';
  tmp_ivl_27825 <= '0';
  tmp_ivl_27837 <= '0';
  tmp_ivl_27844 <= '0';
  tmp_ivl_27860 <= '0';
  tmp_ivl_27867 <= '0';
  tmp_ivl_27879 <= '0';
  tmp_ivl_27888 <= '0';
  tmp_ivl_27902 <= '0';
  tmp_ivl_27913 <= '0';
  tmp_ivl_27925 <= '0';
  tmp_ivl_2793 <= '0';
  tmp_ivl_27932 <= '0';
  tmp_ivl_27944 <= '0';
  tmp_ivl_27951 <= '0';
  tmp_ivl_27967 <= '0';
  tmp_ivl_27974 <= '0';
  tmp_ivl_27986 <= '0';
  tmp_ivl_27995 <= '0';
  tmp_ivl_28009 <= '0';
  tmp_ivl_28020 <= '0';
  tmp_ivl_28032 <= '0';
  tmp_ivl_28039 <= '0';
  tmp_ivl_2804 <= '0';
  tmp_ivl_28051 <= '0';
  tmp_ivl_28058 <= '0';
  tmp_ivl_28074 <= '0';
  tmp_ivl_28081 <= '0';
  tmp_ivl_28093 <= '0';
  tmp_ivl_281 <= '0';
  tmp_ivl_28102 <= '0';
  tmp_ivl_28116 <= '0';
  tmp_ivl_28127 <= '0';
  tmp_ivl_28139 <= '0';
  tmp_ivl_28146 <= '0';
  tmp_ivl_28158 <= '0';
  tmp_ivl_28165 <= '0';
  tmp_ivl_28181 <= '0';
  tmp_ivl_28188 <= '0';
  tmp_ivl_28200 <= '0';
  tmp_ivl_28209 <= '0';
  tmp_ivl_2822 <= '0';
  tmp_ivl_28223 <= '0';
  tmp_ivl_28234 <= '0';
  tmp_ivl_28246 <= '0';
  tmp_ivl_28253 <= '0';
  tmp_ivl_28265 <= '0';
  tmp_ivl_28272 <= '0';
  tmp_ivl_28288 <= '0';
  tmp_ivl_28295 <= '0';
  tmp_ivl_28307 <= '0';
  tmp_ivl_28316 <= '0';
  tmp_ivl_2833 <= '0';
  tmp_ivl_28330 <= '0';
  tmp_ivl_28341 <= '0';
  tmp_ivl_28353 <= '0';
  tmp_ivl_28360 <= '0';
  tmp_ivl_28372 <= '0';
  tmp_ivl_28379 <= '0';
  tmp_ivl_28395 <= '0';
  tmp_ivl_28404 <= '0';
  tmp_ivl_28418 <= '0';
  tmp_ivl_28429 <= '0';
  tmp_ivl_28441 <= '0';
  tmp_ivl_28448 <= '0';
  tmp_ivl_28460 <= '0';
  tmp_ivl_28467 <= '0';
  tmp_ivl_28479 <= '0';
  tmp_ivl_28486 <= '0';
  tmp_ivl_28502 <= '0';
  tmp_ivl_2851 <= '0';
  tmp_ivl_28511 <= '0';
  tmp_ivl_28525 <= '0';
  tmp_ivl_28536 <= '0';
  tmp_ivl_28548 <= '0';
  tmp_ivl_28555 <= '0';
  tmp_ivl_28567 <= '0';
  tmp_ivl_28574 <= '0';
  tmp_ivl_28586 <= '0';
  tmp_ivl_28593 <= '0';
  tmp_ivl_28609 <= '0';
  tmp_ivl_28616 <= '0';
  tmp_ivl_2862 <= '0';
  tmp_ivl_28628 <= '0';
  tmp_ivl_28637 <= '0';
  tmp_ivl_28651 <= '0';
  tmp_ivl_28662 <= '0';
  tmp_ivl_28674 <= '0';
  tmp_ivl_28681 <= '0';
  tmp_ivl_28693 <= '0';
  tmp_ivl_28700 <= '0';
  tmp_ivl_28716 <= '0';
  tmp_ivl_28723 <= '0';
  tmp_ivl_28735 <= '0';
  tmp_ivl_28744 <= '0';
  tmp_ivl_28758 <= '0';
  tmp_ivl_28769 <= '0';
  tmp_ivl_28781 <= '0';
  tmp_ivl_28788 <= '0';
  tmp_ivl_2880 <= '0';
  tmp_ivl_28800 <= '0';
  tmp_ivl_28807 <= '0';
  tmp_ivl_28823 <= '0';
  tmp_ivl_28832 <= '0';
  tmp_ivl_28846 <= '0';
  tmp_ivl_28857 <= '0';
  tmp_ivl_28869 <= '0';
  tmp_ivl_28876 <= '0';
  tmp_ivl_28888 <= '0';
  tmp_ivl_28895 <= '0';
  tmp_ivl_28907 <= '0';
  tmp_ivl_2891 <= '0';
  tmp_ivl_28914 <= '0';
  tmp_ivl_28930 <= '0';
  tmp_ivl_28937 <= '0';
  tmp_ivl_28949 <= '0';
  tmp_ivl_28958 <= '0';
  tmp_ivl_28972 <= '0';
  tmp_ivl_28983 <= '0';
  tmp_ivl_28995 <= '0';
  tmp_ivl_29002 <= '0';
  tmp_ivl_29014 <= '0';
  tmp_ivl_29021 <= '0';
  tmp_ivl_29037 <= '0';
  tmp_ivl_29046 <= '0';
  tmp_ivl_29060 <= '0';
  tmp_ivl_29071 <= '0';
  tmp_ivl_29083 <= '0';
  tmp_ivl_2909 <= '0';
  tmp_ivl_29090 <= '0';
  tmp_ivl_29102 <= '0';
  tmp_ivl_29109 <= '0';
  tmp_ivl_29121 <= '0';
  tmp_ivl_29128 <= '0';
  tmp_ivl_29144 <= '0';
  tmp_ivl_29153 <= '0';
  tmp_ivl_29167 <= '0';
  tmp_ivl_29178 <= '0';
  tmp_ivl_29190 <= '0';
  tmp_ivl_29197 <= '0';
  tmp_ivl_2920 <= '0';
  tmp_ivl_29209 <= '0';
  tmp_ivl_29216 <= '0';
  tmp_ivl_29228 <= '0';
  tmp_ivl_29235 <= '0';
  tmp_ivl_29251 <= '0';
  tmp_ivl_29258 <= '0';
  tmp_ivl_29270 <= '0';
  tmp_ivl_29279 <= '0';
  tmp_ivl_29293 <= '0';
  tmp_ivl_29304 <= '0';
  tmp_ivl_29316 <= '0';
  tmp_ivl_29323 <= '0';
  tmp_ivl_29335 <= '0';
  tmp_ivl_29342 <= '0';
  tmp_ivl_29358 <= '0';
  tmp_ivl_29365 <= '0';
  tmp_ivl_29377 <= '0';
  tmp_ivl_2938 <= '0';
  tmp_ivl_29386 <= '0';
  tmp_ivl_29400 <= '0';
  tmp_ivl_29411 <= '0';
  tmp_ivl_29423 <= '0';
  tmp_ivl_29430 <= '0';
  tmp_ivl_29442 <= '0';
  tmp_ivl_29449 <= '0';
  tmp_ivl_29465 <= '0';
  tmp_ivl_29474 <= '0';
  tmp_ivl_29488 <= '0';
  tmp_ivl_2949 <= '0';
  tmp_ivl_29499 <= '0';
  tmp_ivl_29511 <= '0';
  tmp_ivl_29518 <= '0';
  tmp_ivl_29530 <= '0';
  tmp_ivl_29537 <= '0';
  tmp_ivl_29549 <= '0';
  tmp_ivl_29556 <= '0';
  tmp_ivl_29572 <= '0';
  tmp_ivl_29581 <= '0';
  tmp_ivl_29595 <= '0';
  tmp_ivl_29606 <= '0';
  tmp_ivl_29618 <= '0';
  tmp_ivl_29625 <= '0';
  tmp_ivl_29637 <= '0';
  tmp_ivl_29644 <= '0';
  tmp_ivl_29656 <= '0';
  tmp_ivl_29663 <= '0';
  tmp_ivl_2967 <= '0';
  tmp_ivl_29679 <= '0';
  tmp_ivl_29686 <= '0';
  tmp_ivl_29698 <= '0';
  tmp_ivl_29707 <= '0';
  tmp_ivl_29721 <= '0';
  tmp_ivl_29732 <= '0';
  tmp_ivl_29744 <= '0';
  tmp_ivl_29751 <= '0';
  tmp_ivl_29763 <= '0';
  tmp_ivl_29770 <= '0';
  tmp_ivl_2978 <= '0';
  tmp_ivl_29786 <= '0';
  tmp_ivl_29795 <= '0';
  tmp_ivl_29809 <= '0';
  tmp_ivl_29820 <= '0';
  tmp_ivl_29832 <= '0';
  tmp_ivl_29839 <= '0';
  tmp_ivl_29851 <= '0';
  tmp_ivl_29858 <= '0';
  tmp_ivl_29870 <= '0';
  tmp_ivl_29877 <= '0';
  tmp_ivl_29893 <= '0';
  tmp_ivl_299 <= '0';
  tmp_ivl_29902 <= '0';
  tmp_ivl_29916 <= '0';
  tmp_ivl_29927 <= '0';
  tmp_ivl_29939 <= '0';
  tmp_ivl_29946 <= '0';
  tmp_ivl_29958 <= '0';
  tmp_ivl_2996 <= '0';
  tmp_ivl_29965 <= '0';
  tmp_ivl_29977 <= '0';
  tmp_ivl_29984 <= '0';
  tmp_ivl_30000 <= '0';
  tmp_ivl_30009 <= '0';
  tmp_ivl_30023 <= '0';
  tmp_ivl_30034 <= '0';
  tmp_ivl_30046 <= '0';
  tmp_ivl_30053 <= '0';
  tmp_ivl_30065 <= '0';
  tmp_ivl_3007 <= '0';
  tmp_ivl_30072 <= '0';
  tmp_ivl_30084 <= '0';
  tmp_ivl_30091 <= '0';
  tmp_ivl_30107 <= '0';
  tmp_ivl_30116 <= '0';
  tmp_ivl_30130 <= '0';
  tmp_ivl_30141 <= '0';
  tmp_ivl_30153 <= '0';
  tmp_ivl_30160 <= '0';
  tmp_ivl_30172 <= '0';
  tmp_ivl_30179 <= '0';
  tmp_ivl_30191 <= '0';
  tmp_ivl_30198 <= '0';
  tmp_ivl_30214 <= '0';
  tmp_ivl_30223 <= '0';
  tmp_ivl_30237 <= '0';
  tmp_ivl_30248 <= '0';
  tmp_ivl_3025 <= '0';
  tmp_ivl_30260 <= '0';
  tmp_ivl_30267 <= '0';
  tmp_ivl_30279 <= '0';
  tmp_ivl_30286 <= '0';
  tmp_ivl_30298 <= '0';
  tmp_ivl_30305 <= '0';
  tmp_ivl_30323 <= '0';
  tmp_ivl_30330 <= '0';
  tmp_ivl_30337 <= '0';
  tmp_ivl_30346 <= '0';
  tmp_ivl_30353 <= '0';
  tmp_ivl_3036 <= '0';
  tmp_ivl_30365 <= '0';
  tmp_ivl_30374 <= '0';
  tmp_ivl_30386 <= '0';
  tmp_ivl_30397 <= '0';
  tmp_ivl_30409 <= '0';
  tmp_ivl_30416 <= '0';
  tmp_ivl_30428 <= '0';
  tmp_ivl_30435 <= '0';
  tmp_ivl_30451 <= '0';
  tmp_ivl_30458 <= '0';
  tmp_ivl_30470 <= '0';
  tmp_ivl_30477 <= '0';
  tmp_ivl_30493 <= '0';
  tmp_ivl_30502 <= '0';
  tmp_ivl_30516 <= '0';
  tmp_ivl_30527 <= '0';
  tmp_ivl_30539 <= '0';
  tmp_ivl_3054 <= '0';
  tmp_ivl_30546 <= '0';
  tmp_ivl_30558 <= '0';
  tmp_ivl_30565 <= '0';
  tmp_ivl_30577 <= '0';
  tmp_ivl_30584 <= '0';
  tmp_ivl_30600 <= '0';
  tmp_ivl_30609 <= '0';
  tmp_ivl_30623 <= '0';
  tmp_ivl_30634 <= '0';
  tmp_ivl_30646 <= '0';
  tmp_ivl_3065 <= '0';
  tmp_ivl_30653 <= '0';
  tmp_ivl_30665 <= '0';
  tmp_ivl_30672 <= '0';
  tmp_ivl_30684 <= '0';
  tmp_ivl_30691 <= '0';
  tmp_ivl_30707 <= '0';
  tmp_ivl_30716 <= '0';
  tmp_ivl_30728 <= '0';
  tmp_ivl_30737 <= '0';
  tmp_ivl_30749 <= '0';
  tmp_ivl_30760 <= '0';
  tmp_ivl_30772 <= '0';
  tmp_ivl_30779 <= '0';
  tmp_ivl_30791 <= '0';
  tmp_ivl_30798 <= '0';
  tmp_ivl_30814 <= '0';
  tmp_ivl_30821 <= '0';
  tmp_ivl_3083 <= '0';
  tmp_ivl_30833 <= '0';
  tmp_ivl_30840 <= '0';
  tmp_ivl_30858 <= '0';
  tmp_ivl_30865 <= '0';
  tmp_ivl_30877 <= '0';
  tmp_ivl_30886 <= '0';
  tmp_ivl_30898 <= '0';
  tmp_ivl_30905 <= '0';
  tmp_ivl_30917 <= '0';
  tmp_ivl_30924 <= '0';
  tmp_ivl_3094 <= '0';
  tmp_ivl_30940 <= '0';
  tmp_ivl_30947 <= '0';
  tmp_ivl_30961 <= '0';
  tmp_ivl_30972 <= '0';
  tmp_ivl_30984 <= '0';
  tmp_ivl_30991 <= '0';
  tmp_ivl_310 <= '0';
  tmp_ivl_31003 <= '0';
  tmp_ivl_31010 <= '0';
  tmp_ivl_31026 <= '0';
  tmp_ivl_31033 <= '0';
  tmp_ivl_31045 <= '0';
  tmp_ivl_31052 <= '0';
  tmp_ivl_31070 <= '0';
  tmp_ivl_31077 <= '0';
  tmp_ivl_31084 <= '0';
  tmp_ivl_31091 <= '0';
  tmp_ivl_31098 <= '0';
  tmp_ivl_31110 <= '0';
  tmp_ivl_31119 <= '0';
  tmp_ivl_3112 <= '0';
  tmp_ivl_31135 <= '0';
  tmp_ivl_31142 <= '0';
  tmp_ivl_31154 <= '0';
  tmp_ivl_31161 <= '0';
  tmp_ivl_31173 <= '0';
  tmp_ivl_31180 <= '0';
  tmp_ivl_31196 <= '0';
  tmp_ivl_31203 <= '0';
  tmp_ivl_31215 <= '0';
  tmp_ivl_31222 <= '0';
  tmp_ivl_3123 <= '0';
  tmp_ivl_31238 <= '0';
  tmp_ivl_31245 <= '0';
  tmp_ivl_31257 <= '0';
  tmp_ivl_31264 <= '0';
  tmp_ivl_31282 <= '0';
  tmp_ivl_31289 <= '0';
  tmp_ivl_31303 <= '0';
  tmp_ivl_31314 <= '0';
  tmp_ivl_31326 <= '0';
  tmp_ivl_31333 <= '0';
  tmp_ivl_31345 <= '0';
  tmp_ivl_31352 <= '0';
  tmp_ivl_31364 <= '0';
  tmp_ivl_31371 <= '0';
  tmp_ivl_31387 <= '0';
  tmp_ivl_31394 <= '0';
  tmp_ivl_31406 <= '0';
  tmp_ivl_3141 <= '0';
  tmp_ivl_31413 <= '0';
  tmp_ivl_31429 <= '0';
  tmp_ivl_31436 <= '0';
  tmp_ivl_31448 <= '0';
  tmp_ivl_31455 <= '0';
  tmp_ivl_31473 <= '0';
  tmp_ivl_31480 <= '0';
  tmp_ivl_31492 <= '0';
  tmp_ivl_31499 <= '0';
  tmp_ivl_31511 <= '0';
  tmp_ivl_31518 <= '0';
  tmp_ivl_3152 <= '0';
  tmp_ivl_31534 <= '0';
  tmp_ivl_31541 <= '0';
  tmp_ivl_31553 <= '0';
  tmp_ivl_31560 <= '0';
  tmp_ivl_31576 <= '0';
  tmp_ivl_31585 <= '0';
  tmp_ivl_31597 <= '0';
  tmp_ivl_31604 <= '0';
  tmp_ivl_31616 <= '0';
  tmp_ivl_31625 <= '0';
  tmp_ivl_31637 <= '0';
  tmp_ivl_31644 <= '0';
  tmp_ivl_31662 <= '0';
  tmp_ivl_31673 <= '0';
  tmp_ivl_31685 <= '0';
  tmp_ivl_31692 <= '0';
  tmp_ivl_3170 <= '0';
  tmp_ivl_31704 <= '0';
  tmp_ivl_31711 <= '0';
  tmp_ivl_31723 <= '0';
  tmp_ivl_31730 <= '0';
  tmp_ivl_31746 <= '0';
  tmp_ivl_31753 <= '0';
  tmp_ivl_31765 <= '0';
  tmp_ivl_31772 <= '0';
  tmp_ivl_31788 <= '0';
  tmp_ivl_31795 <= '0';
  tmp_ivl_31807 <= '0';
  tmp_ivl_3181 <= '0';
  tmp_ivl_31814 <= '0';
  tmp_ivl_31830 <= '0';
  tmp_ivl_31837 <= '0';
  tmp_ivl_31851 <= '0';
  tmp_ivl_31858 <= '0';
  tmp_ivl_31865 <= '0';
  tmp_ivl_31874 <= '0';
  tmp_ivl_31881 <= '0';
  tmp_ivl_31893 <= '0';
  tmp_ivl_31900 <= '0';
  tmp_ivl_31916 <= '0';
  tmp_ivl_31923 <= '0';
  tmp_ivl_31935 <= '0';
  tmp_ivl_31942 <= '0';
  tmp_ivl_31949 <= '0';
  tmp_ivl_31958 <= '0';
  tmp_ivl_31965 <= '0';
  tmp_ivl_31981 <= '0';
  tmp_ivl_31988 <= '0';
  tmp_ivl_3199 <= '0';
  tmp_ivl_32000 <= '0';
  tmp_ivl_32007 <= '0';
  tmp_ivl_32023 <= '0';
  tmp_ivl_32030 <= '0';
  tmp_ivl_32042 <= '0';
  tmp_ivl_32049 <= '0';
  tmp_ivl_32065 <= '0';
  tmp_ivl_32072 <= '0';
  tmp_ivl_32084 <= '0';
  tmp_ivl_32091 <= '0';
  tmp_ivl_3210 <= '0';
  tmp_ivl_32107 <= '0';
  tmp_ivl_32114 <= '0';
  tmp_ivl_32126 <= '0';
  tmp_ivl_32133 <= '0';
  tmp_ivl_32149 <= '0';
  tmp_ivl_32156 <= '0';
  tmp_ivl_32168 <= '0';
  tmp_ivl_32175 <= '0';
  tmp_ivl_32191 <= '0';
  tmp_ivl_32198 <= '0';
  tmp_ivl_32210 <= '0';
  tmp_ivl_32217 <= '0';
  tmp_ivl_32233 <= '0';
  tmp_ivl_32240 <= '0';
  tmp_ivl_32252 <= '0';
  tmp_ivl_32259 <= '0';
  tmp_ivl_32275 <= '0';
  tmp_ivl_3228 <= '0';
  tmp_ivl_32282 <= '0';
  tmp_ivl_32294 <= '0';
  tmp_ivl_32301 <= '0';
  tmp_ivl_32317 <= '0';
  tmp_ivl_32324 <= '0';
  tmp_ivl_32336 <= '0';
  tmp_ivl_32343 <= '0';
  tmp_ivl_32359 <= '0';
  tmp_ivl_32366 <= '0';
  tmp_ivl_32378 <= '0';
  tmp_ivl_32385 <= '0';
  tmp_ivl_3239 <= '0';
  tmp_ivl_32401 <= '0';
  tmp_ivl_32408 <= '0';
  tmp_ivl_32420 <= '0';
  tmp_ivl_32427 <= '0';
  tmp_ivl_32443 <= '0';
  tmp_ivl_32450 <= '0';
  tmp_ivl_32462 <= '0';
  tmp_ivl_32469 <= '0';
  tmp_ivl_32485 <= '0';
  tmp_ivl_32492 <= '0';
  tmp_ivl_32504 <= '0';
  tmp_ivl_32511 <= '0';
  tmp_ivl_32527 <= '0';
  tmp_ivl_32534 <= '0';
  tmp_ivl_32546 <= '0';
  tmp_ivl_32553 <= '0';
  tmp_ivl_32569 <= '0';
  tmp_ivl_3257 <= '0';
  tmp_ivl_32576 <= '0';
  tmp_ivl_32588 <= '0';
  tmp_ivl_32595 <= '0';
  tmp_ivl_32611 <= '0';
  tmp_ivl_32618 <= '0';
  tmp_ivl_32630 <= '0';
  tmp_ivl_32637 <= '0';
  tmp_ivl_32653 <= '0';
  tmp_ivl_32660 <= '0';
  tmp_ivl_32672 <= '0';
  tmp_ivl_32679 <= '0';
  tmp_ivl_3268 <= '0';
  tmp_ivl_32695 <= '0';
  tmp_ivl_32702 <= '0';
  tmp_ivl_32714 <= '0';
  tmp_ivl_32721 <= '0';
  tmp_ivl_32737 <= '0';
  tmp_ivl_32744 <= '0';
  tmp_ivl_32756 <= '0';
  tmp_ivl_32763 <= '0';
  tmp_ivl_32779 <= '0';
  tmp_ivl_32786 <= '0';
  tmp_ivl_32798 <= '0';
  tmp_ivl_328 <= '0';
  tmp_ivl_32805 <= '0';
  tmp_ivl_32821 <= '0';
  tmp_ivl_32828 <= '0';
  tmp_ivl_32840 <= '0';
  tmp_ivl_32847 <= '0';
  tmp_ivl_3286 <= '0';
  tmp_ivl_32863 <= '0';
  tmp_ivl_32870 <= '0';
  tmp_ivl_32882 <= '0';
  tmp_ivl_32889 <= '0';
  tmp_ivl_32905 <= '0';
  tmp_ivl_32912 <= '0';
  tmp_ivl_32924 <= '0';
  tmp_ivl_32931 <= '0';
  tmp_ivl_32947 <= '0';
  tmp_ivl_32954 <= '0';
  tmp_ivl_32966 <= '0';
  tmp_ivl_3297 <= '0';
  tmp_ivl_32973 <= '0';
  tmp_ivl_32989 <= '0';
  tmp_ivl_32996 <= '0';
  tmp_ivl_33008 <= '0';
  tmp_ivl_33015 <= '0';
  tmp_ivl_33031 <= '0';
  tmp_ivl_33038 <= '0';
  tmp_ivl_33050 <= '0';
  tmp_ivl_33057 <= '0';
  tmp_ivl_33073 <= '0';
  tmp_ivl_33080 <= '0';
  tmp_ivl_33092 <= '0';
  tmp_ivl_33099 <= '0';
  tmp_ivl_33115 <= '0';
  tmp_ivl_33122 <= '0';
  tmp_ivl_33134 <= '0';
  tmp_ivl_33141 <= '0';
  tmp_ivl_3315 <= '0';
  tmp_ivl_33157 <= '0';
  tmp_ivl_33164 <= '0';
  tmp_ivl_33176 <= '0';
  tmp_ivl_33183 <= '0';
  tmp_ivl_33199 <= '0';
  tmp_ivl_33206 <= '0';
  tmp_ivl_33218 <= '0';
  tmp_ivl_33225 <= '0';
  tmp_ivl_33241 <= '0';
  tmp_ivl_33248 <= '0';
  tmp_ivl_3326 <= '0';
  tmp_ivl_33260 <= '0';
  tmp_ivl_33267 <= '0';
  tmp_ivl_33283 <= '0';
  tmp_ivl_33290 <= '0';
  tmp_ivl_33302 <= '0';
  tmp_ivl_33309 <= '0';
  tmp_ivl_33325 <= '0';
  tmp_ivl_33332 <= '0';
  tmp_ivl_33344 <= '0';
  tmp_ivl_33351 <= '0';
  tmp_ivl_33367 <= '0';
  tmp_ivl_33374 <= '0';
  tmp_ivl_33386 <= '0';
  tmp_ivl_33393 <= '0';
  tmp_ivl_33409 <= '0';
  tmp_ivl_33416 <= '0';
  tmp_ivl_33428 <= '0';
  tmp_ivl_33435 <= '0';
  tmp_ivl_3344 <= '0';
  tmp_ivl_33451 <= '0';
  tmp_ivl_33458 <= '0';
  tmp_ivl_33470 <= '0';
  tmp_ivl_33477 <= '0';
  tmp_ivl_33493 <= '0';
  tmp_ivl_33500 <= '0';
  tmp_ivl_33512 <= '0';
  tmp_ivl_33519 <= '0';
  tmp_ivl_33535 <= '0';
  tmp_ivl_33542 <= '0';
  tmp_ivl_3355 <= '0';
  tmp_ivl_33554 <= '0';
  tmp_ivl_33561 <= '0';
  tmp_ivl_33577 <= '0';
  tmp_ivl_33584 <= '0';
  tmp_ivl_33596 <= '0';
  tmp_ivl_33603 <= '0';
  tmp_ivl_33619 <= '0';
  tmp_ivl_33626 <= '0';
  tmp_ivl_33638 <= '0';
  tmp_ivl_33645 <= '0';
  tmp_ivl_33661 <= '0';
  tmp_ivl_33668 <= '0';
  tmp_ivl_33680 <= '0';
  tmp_ivl_33687 <= '0';
  tmp_ivl_33703 <= '0';
  tmp_ivl_33710 <= '0';
  tmp_ivl_33722 <= '0';
  tmp_ivl_33729 <= '0';
  tmp_ivl_3373 <= '0';
  tmp_ivl_33745 <= '0';
  tmp_ivl_33752 <= '0';
  tmp_ivl_33764 <= '0';
  tmp_ivl_33771 <= '0';
  tmp_ivl_33787 <= '0';
  tmp_ivl_33794 <= '0';
  tmp_ivl_33806 <= '0';
  tmp_ivl_33813 <= '0';
  tmp_ivl_33829 <= '0';
  tmp_ivl_33836 <= '0';
  tmp_ivl_3384 <= '0';
  tmp_ivl_33848 <= '0';
  tmp_ivl_33855 <= '0';
  tmp_ivl_33871 <= '0';
  tmp_ivl_33878 <= '0';
  tmp_ivl_33890 <= '0';
  tmp_ivl_33897 <= '0';
  tmp_ivl_339 <= '0';
  tmp_ivl_33913 <= '0';
  tmp_ivl_33920 <= '0';
  tmp_ivl_33932 <= '0';
  tmp_ivl_33939 <= '0';
  tmp_ivl_33955 <= '0';
  tmp_ivl_33962 <= '0';
  tmp_ivl_33974 <= '0';
  tmp_ivl_33981 <= '0';
  tmp_ivl_33997 <= '0';
  tmp_ivl_34004 <= '0';
  tmp_ivl_34016 <= '0';
  tmp_ivl_3402 <= '0';
  tmp_ivl_34023 <= '0';
  tmp_ivl_34039 <= '0';
  tmp_ivl_34046 <= '0';
  tmp_ivl_34058 <= '0';
  tmp_ivl_34065 <= '0';
  tmp_ivl_34081 <= '0';
  tmp_ivl_34088 <= '0';
  tmp_ivl_34100 <= '0';
  tmp_ivl_34107 <= '0';
  tmp_ivl_34123 <= '0';
  tmp_ivl_3413 <= '0';
  tmp_ivl_34130 <= '0';
  tmp_ivl_34137 <= '0';
  tmp_ivl_34144 <= '0';
  tmp_ivl_34151 <= '0';
  tmp_ivl_34163 <= '0';
  tmp_ivl_34170 <= '0';
  tmp_ivl_34186 <= '0';
  tmp_ivl_34195 <= '0';
  tmp_ivl_34207 <= '0';
  tmp_ivl_34214 <= '0';
  tmp_ivl_34226 <= '0';
  tmp_ivl_34233 <= '0';
  tmp_ivl_34249 <= '0';
  tmp_ivl_34256 <= '0';
  tmp_ivl_34268 <= '0';
  tmp_ivl_34275 <= '0';
  tmp_ivl_34291 <= '0';
  tmp_ivl_34298 <= '0';
  tmp_ivl_3431 <= '0';
  tmp_ivl_34310 <= '0';
  tmp_ivl_34317 <= '0';
  tmp_ivl_34333 <= '0';
  tmp_ivl_34340 <= '0';
  tmp_ivl_34352 <= '0';
  tmp_ivl_34359 <= '0';
  tmp_ivl_34375 <= '0';
  tmp_ivl_34382 <= '0';
  tmp_ivl_34394 <= '0';
  tmp_ivl_34401 <= '0';
  tmp_ivl_34417 <= '0';
  tmp_ivl_3442 <= '0';
  tmp_ivl_34424 <= '0';
  tmp_ivl_34436 <= '0';
  tmp_ivl_34443 <= '0';
  tmp_ivl_34461 <= '0';
  tmp_ivl_34472 <= '0';
  tmp_ivl_34484 <= '0';
  tmp_ivl_34491 <= '0';
  tmp_ivl_34503 <= '0';
  tmp_ivl_34510 <= '0';
  tmp_ivl_34522 <= '0';
  tmp_ivl_34529 <= '0';
  tmp_ivl_34545 <= '0';
  tmp_ivl_34552 <= '0';
  tmp_ivl_34564 <= '0';
  tmp_ivl_34571 <= '0';
  tmp_ivl_34587 <= '0';
  tmp_ivl_34594 <= '0';
  tmp_ivl_3460 <= '0';
  tmp_ivl_34606 <= '0';
  tmp_ivl_34613 <= '0';
  tmp_ivl_34631 <= '0';
  tmp_ivl_34642 <= '0';
  tmp_ivl_34654 <= '0';
  tmp_ivl_34661 <= '0';
  tmp_ivl_34673 <= '0';
  tmp_ivl_34680 <= '0';
  tmp_ivl_34692 <= '0';
  tmp_ivl_34699 <= '0';
  tmp_ivl_3471 <= '0';
  tmp_ivl_34715 <= '0';
  tmp_ivl_34722 <= '0';
  tmp_ivl_34734 <= '0';
  tmp_ivl_34741 <= '0';
  tmp_ivl_34757 <= '0';
  tmp_ivl_34764 <= '0';
  tmp_ivl_34776 <= '0';
  tmp_ivl_34783 <= '0';
  tmp_ivl_34801 <= '0';
  tmp_ivl_34812 <= '0';
  tmp_ivl_34824 <= '0';
  tmp_ivl_34831 <= '0';
  tmp_ivl_34843 <= '0';
  tmp_ivl_34850 <= '0';
  tmp_ivl_34862 <= '0';
  tmp_ivl_34869 <= '0';
  tmp_ivl_34885 <= '0';
  tmp_ivl_3489 <= '0';
  tmp_ivl_34892 <= '0';
  tmp_ivl_34904 <= '0';
  tmp_ivl_34911 <= '0';
  tmp_ivl_34927 <= '0';
  tmp_ivl_34934 <= '0';
  tmp_ivl_34946 <= '0';
  tmp_ivl_34953 <= '0';
  tmp_ivl_34971 <= '0';
  tmp_ivl_34982 <= '0';
  tmp_ivl_34994 <= '0';
  tmp_ivl_3500 <= '0';
  tmp_ivl_35001 <= '0';
  tmp_ivl_35013 <= '0';
  tmp_ivl_35020 <= '0';
  tmp_ivl_35032 <= '0';
  tmp_ivl_35039 <= '0';
  tmp_ivl_35055 <= '0';
  tmp_ivl_35062 <= '0';
  tmp_ivl_35074 <= '0';
  tmp_ivl_35081 <= '0';
  tmp_ivl_35097 <= '0';
  tmp_ivl_35104 <= '0';
  tmp_ivl_35116 <= '0';
  tmp_ivl_35123 <= '0';
  tmp_ivl_35141 <= '0';
  tmp_ivl_35148 <= '0';
  tmp_ivl_35155 <= "00";
  tmp_ivl_35169 <= '0';
  tmp_ivl_35176 <= '0';
  tmp_ivl_3518 <= '0';
  tmp_ivl_35183 <= "00";
  tmp_ivl_35197 <= '0';
  tmp_ivl_35204 <= '0';
  tmp_ivl_35211 <= "00";
  tmp_ivl_35225 <= '0';
  tmp_ivl_35232 <= '0';
  tmp_ivl_35239 <= "00";
  tmp_ivl_35253 <= '0';
  tmp_ivl_35260 <= '0';
  tmp_ivl_35267 <= "00";
  tmp_ivl_35281 <= '0';
  tmp_ivl_35288 <= '0';
  tmp_ivl_3529 <= '0';
  tmp_ivl_35295 <= "00";
  tmp_ivl_35309 <= '0';
  tmp_ivl_35316 <= '0';
  tmp_ivl_35323 <= "00";
  tmp_ivl_35337 <= '0';
  tmp_ivl_35344 <= '0';
  tmp_ivl_35351 <= "00";
  tmp_ivl_35365 <= '0';
  tmp_ivl_35372 <= '0';
  tmp_ivl_35379 <= "00";
  tmp_ivl_35393 <= '0';
  tmp_ivl_35400 <= '0';
  tmp_ivl_35407 <= "00";
  tmp_ivl_35421 <= '0';
  tmp_ivl_35428 <= '0';
  tmp_ivl_35435 <= "00";
  tmp_ivl_35451 <= '0';
  tmp_ivl_35458 <= '0';
  tmp_ivl_35465 <= "00";
  tmp_ivl_3547 <= '0';
  tmp_ivl_35479 <= '0';
  tmp_ivl_35486 <= '0';
  tmp_ivl_35493 <= "00";
  tmp_ivl_35507 <= '0';
  tmp_ivl_35514 <= '0';
  tmp_ivl_35521 <= "00";
  tmp_ivl_35535 <= '0';
  tmp_ivl_35542 <= '0';
  tmp_ivl_35549 <= "00";
  tmp_ivl_35563 <= '0';
  tmp_ivl_35570 <= '0';
  tmp_ivl_35577 <= "00";
  tmp_ivl_3558 <= '0';
  tmp_ivl_35591 <= '0';
  tmp_ivl_35598 <= '0';
  tmp_ivl_35605 <= "00";
  tmp_ivl_35619 <= '0';
  tmp_ivl_35626 <= '0';
  tmp_ivl_35633 <= "00";
  tmp_ivl_35647 <= '0';
  tmp_ivl_35654 <= '0';
  tmp_ivl_35661 <= "00";
  tmp_ivl_35675 <= '0';
  tmp_ivl_35682 <= '0';
  tmp_ivl_35689 <= "00";
  tmp_ivl_357 <= '0';
  tmp_ivl_35703 <= '0';
  tmp_ivl_35710 <= '0';
  tmp_ivl_35717 <= "00";
  tmp_ivl_35731 <= '0';
  tmp_ivl_35738 <= '0';
  tmp_ivl_35745 <= "00";
  tmp_ivl_35759 <= '0';
  tmp_ivl_3576 <= '0';
  tmp_ivl_35766 <= '0';
  tmp_ivl_35773 <= "00";
  tmp_ivl_35787 <= '0';
  tmp_ivl_35794 <= '0';
  tmp_ivl_35801 <= "00";
  tmp_ivl_35815 <= '0';
  tmp_ivl_35822 <= '0';
  tmp_ivl_35829 <= "00";
  tmp_ivl_35843 <= '0';
  tmp_ivl_35850 <= '0';
  tmp_ivl_35857 <= "00";
  tmp_ivl_3587 <= '0';
  tmp_ivl_35871 <= '0';
  tmp_ivl_35878 <= '0';
  tmp_ivl_35885 <= "00";
  tmp_ivl_35899 <= '0';
  tmp_ivl_35906 <= '0';
  tmp_ivl_35913 <= "00";
  tmp_ivl_35927 <= '0';
  tmp_ivl_35934 <= '0';
  tmp_ivl_35941 <= "00";
  tmp_ivl_35955 <= '0';
  tmp_ivl_35962 <= '0';
  tmp_ivl_35969 <= "00";
  tmp_ivl_35983 <= '0';
  tmp_ivl_35990 <= '0';
  tmp_ivl_35997 <= "00";
  tmp_ivl_36011 <= '0';
  tmp_ivl_36018 <= '0';
  tmp_ivl_36025 <= "00";
  tmp_ivl_36039 <= '0';
  tmp_ivl_36046 <= '0';
  tmp_ivl_3605 <= '0';
  tmp_ivl_36053 <= "00";
  tmp_ivl_36067 <= '0';
  tmp_ivl_36074 <= '0';
  tmp_ivl_36081 <= "00";
  tmp_ivl_36095 <= '0';
  tmp_ivl_36102 <= '0';
  tmp_ivl_36109 <= "00";
  tmp_ivl_36123 <= '0';
  tmp_ivl_36130 <= '0';
  tmp_ivl_36137 <= "00";
  tmp_ivl_36151 <= '0';
  tmp_ivl_36158 <= '0';
  tmp_ivl_3616 <= '0';
  tmp_ivl_36165 <= "00";
  tmp_ivl_36179 <= '0';
  tmp_ivl_36186 <= '0';
  tmp_ivl_36193 <= "00";
  tmp_ivl_36207 <= '0';
  tmp_ivl_36214 <= '0';
  tmp_ivl_36221 <= "00";
  tmp_ivl_36235 <= '0';
  tmp_ivl_36242 <= '0';
  tmp_ivl_36249 <= "00";
  tmp_ivl_36263 <= '0';
  tmp_ivl_36270 <= '0';
  tmp_ivl_36277 <= "00";
  tmp_ivl_36291 <= '0';
  tmp_ivl_36298 <= '0';
  tmp_ivl_36305 <= "00";
  tmp_ivl_36319 <= '0';
  tmp_ivl_36326 <= '0';
  tmp_ivl_36333 <= "00";
  tmp_ivl_3634 <= '0';
  tmp_ivl_36347 <= '0';
  tmp_ivl_36354 <= '0';
  tmp_ivl_36361 <= "00";
  tmp_ivl_36375 <= '0';
  tmp_ivl_36382 <= '0';
  tmp_ivl_36389 <= "00";
  tmp_ivl_36403 <= '0';
  tmp_ivl_36410 <= '0';
  tmp_ivl_36417 <= "00";
  tmp_ivl_36431 <= '0';
  tmp_ivl_36438 <= '0';
  tmp_ivl_36445 <= "00";
  tmp_ivl_3645 <= '0';
  tmp_ivl_36459 <= '0';
  tmp_ivl_36466 <= '0';
  tmp_ivl_36473 <= "00";
  tmp_ivl_36487 <= '0';
  tmp_ivl_36494 <= '0';
  tmp_ivl_36501 <= "00";
  tmp_ivl_36515 <= '0';
  tmp_ivl_36522 <= '0';
  tmp_ivl_36529 <= "00";
  tmp_ivl_36543 <= '0';
  tmp_ivl_36550 <= '0';
  tmp_ivl_36557 <= "00";
  tmp_ivl_36571 <= '0';
  tmp_ivl_36578 <= '0';
  tmp_ivl_36585 <= "00";
  tmp_ivl_36599 <= '0';
  tmp_ivl_36606 <= '0';
  tmp_ivl_36613 <= "00";
  tmp_ivl_36627 <= '0';
  tmp_ivl_3663 <= '0';
  tmp_ivl_36634 <= '0';
  tmp_ivl_36641 <= "00";
  tmp_ivl_36655 <= '0';
  tmp_ivl_36662 <= '0';
  tmp_ivl_36669 <= "00";
  tmp_ivl_36683 <= '0';
  tmp_ivl_36690 <= '0';
  tmp_ivl_36697 <= "00";
  tmp_ivl_36711 <= '0';
  tmp_ivl_36718 <= '0';
  tmp_ivl_36725 <= "00";
  tmp_ivl_36739 <= '0';
  tmp_ivl_3674 <= '0';
  tmp_ivl_36746 <= '0';
  tmp_ivl_36753 <= "00";
  tmp_ivl_36767 <= '0';
  tmp_ivl_36774 <= '0';
  tmp_ivl_36781 <= "00";
  tmp_ivl_36795 <= '0';
  tmp_ivl_368 <= '0';
  tmp_ivl_36802 <= '0';
  tmp_ivl_36809 <= "00";
  tmp_ivl_36823 <= '0';
  tmp_ivl_36830 <= '0';
  tmp_ivl_36837 <= "00";
  tmp_ivl_36851 <= '0';
  tmp_ivl_36858 <= '0';
  tmp_ivl_36865 <= "00";
  tmp_ivl_36879 <= '0';
  tmp_ivl_36886 <= '0';
  tmp_ivl_36893 <= "00";
  tmp_ivl_36907 <= '0';
  tmp_ivl_36914 <= '0';
  tmp_ivl_3692 <= '0';
  tmp_ivl_36921 <= "00";
  tmp_ivl_36937 <= '0';
  tmp_ivl_36944 <= '0';
  tmp_ivl_36951 <= "00";
  tmp_ivl_36967 <= '0';
  tmp_ivl_36974 <= '0';
  tmp_ivl_36981 <= "00";
  tmp_ivl_36997 <= '0';
  tmp_ivl_37004 <= '0';
  tmp_ivl_37011 <= "00";
  tmp_ivl_37027 <= '0';
  tmp_ivl_3703 <= '0';
  tmp_ivl_37034 <= '0';
  tmp_ivl_37041 <= "00";
  tmp_ivl_37057 <= '0';
  tmp_ivl_37064 <= '0';
  tmp_ivl_37071 <= "00";
  tmp_ivl_37087 <= '0';
  tmp_ivl_37094 <= '0';
  tmp_ivl_37101 <= "00";
  tmp_ivl_37117 <= '0';
  tmp_ivl_37124 <= '0';
  tmp_ivl_37131 <= "00";
  tmp_ivl_37147 <= '0';
  tmp_ivl_37154 <= '0';
  tmp_ivl_37161 <= "00";
  tmp_ivl_37177 <= '0';
  tmp_ivl_37184 <= '0';
  tmp_ivl_37191 <= "00";
  tmp_ivl_37207 <= '0';
  tmp_ivl_3721 <= '0';
  tmp_ivl_37214 <= '0';
  tmp_ivl_37221 <= "00";
  tmp_ivl_37237 <= '0';
  tmp_ivl_37244 <= '0';
  tmp_ivl_37251 <= "00";
  tmp_ivl_37267 <= '0';
  tmp_ivl_37274 <= '0';
  tmp_ivl_37281 <= "00";
  tmp_ivl_37297 <= '0';
  tmp_ivl_37304 <= '0';
  tmp_ivl_37311 <= "00";
  tmp_ivl_3732 <= '0';
  tmp_ivl_37327 <= '0';
  tmp_ivl_37334 <= '0';
  tmp_ivl_37341 <= "00";
  tmp_ivl_37357 <= '0';
  tmp_ivl_37364 <= '0';
  tmp_ivl_37371 <= "00";
  tmp_ivl_37387 <= '0';
  tmp_ivl_37394 <= '0';
  tmp_ivl_37401 <= "00";
  tmp_ivl_37417 <= '0';
  tmp_ivl_37424 <= '0';
  tmp_ivl_37431 <= "00";
  tmp_ivl_37447 <= '0';
  tmp_ivl_37454 <= '0';
  tmp_ivl_37461 <= "00";
  tmp_ivl_37477 <= '0';
  tmp_ivl_3748 <= '0';
  tmp_ivl_37484 <= '0';
  tmp_ivl_37491 <= "00";
  tmp_ivl_37507 <= '0';
  tmp_ivl_37514 <= '0';
  tmp_ivl_37521 <= "00";
  tmp_ivl_37537 <= '0';
  tmp_ivl_37544 <= '0';
  tmp_ivl_37551 <= "00";
  tmp_ivl_37567 <= '0';
  tmp_ivl_37574 <= '0';
  tmp_ivl_37581 <= "00";
  tmp_ivl_3759 <= '0';
  tmp_ivl_37597 <= '0';
  tmp_ivl_37604 <= '0';
  tmp_ivl_37611 <= "00";
  tmp_ivl_37627 <= '0';
  tmp_ivl_37634 <= '0';
  tmp_ivl_37641 <= "00";
  tmp_ivl_37657 <= '0';
  tmp_ivl_37664 <= '0';
  tmp_ivl_37671 <= "00";
  tmp_ivl_37687 <= '0';
  tmp_ivl_37694 <= '0';
  tmp_ivl_37701 <= "00";
  tmp_ivl_37717 <= '0';
  tmp_ivl_37724 <= '0';
  tmp_ivl_37731 <= "00";
  tmp_ivl_37747 <= '0';
  tmp_ivl_3775 <= '0';
  tmp_ivl_37754 <= '0';
  tmp_ivl_37761 <= "00";
  tmp_ivl_37777 <= '0';
  tmp_ivl_37784 <= '0';
  tmp_ivl_37791 <= "00";
  tmp_ivl_37807 <= '0';
  tmp_ivl_37814 <= '0';
  tmp_ivl_37821 <= "00";
  tmp_ivl_37837 <= '0';
  tmp_ivl_37844 <= '0';
  tmp_ivl_37851 <= "00";
  tmp_ivl_3786 <= '0';
  tmp_ivl_37867 <= '0';
  tmp_ivl_37874 <= '0';
  tmp_ivl_37881 <= "00";
  tmp_ivl_37897 <= '0';
  tmp_ivl_37904 <= '0';
  tmp_ivl_37911 <= "00";
  tmp_ivl_37927 <= '0';
  tmp_ivl_37934 <= '0';
  tmp_ivl_37941 <= "00";
  tmp_ivl_37957 <= '0';
  tmp_ivl_37964 <= '0';
  tmp_ivl_37971 <= "00";
  tmp_ivl_37987 <= '0';
  tmp_ivl_37994 <= '0';
  tmp_ivl_38 <= '0';
  tmp_ivl_38001 <= "00";
  tmp_ivl_38017 <= '0';
  tmp_ivl_3802 <= '0';
  tmp_ivl_38024 <= '0';
  tmp_ivl_38031 <= "00";
  tmp_ivl_38047 <= '0';
  tmp_ivl_38054 <= '0';
  tmp_ivl_38061 <= "00";
  tmp_ivl_38077 <= '0';
  tmp_ivl_38084 <= '0';
  tmp_ivl_38091 <= "00";
  tmp_ivl_38107 <= '0';
  tmp_ivl_38114 <= '0';
  tmp_ivl_38121 <= "00";
  tmp_ivl_3813 <= '0';
  tmp_ivl_38137 <= '0';
  tmp_ivl_38144 <= '0';
  tmp_ivl_38151 <= "00";
  tmp_ivl_38167 <= '0';
  tmp_ivl_38174 <= '0';
  tmp_ivl_38181 <= "00";
  tmp_ivl_38197 <= '0';
  tmp_ivl_38204 <= '0';
  tmp_ivl_38211 <= "00";
  tmp_ivl_38227 <= '0';
  tmp_ivl_38234 <= '0';
  tmp_ivl_38241 <= "00";
  tmp_ivl_38257 <= '0';
  tmp_ivl_38264 <= '0';
  tmp_ivl_38271 <= "00";
  tmp_ivl_38287 <= '0';
  tmp_ivl_3829 <= '0';
  tmp_ivl_38294 <= '0';
  tmp_ivl_38301 <= "00";
  tmp_ivl_38317 <= '0';
  tmp_ivl_38324 <= '0';
  tmp_ivl_38331 <= "00";
  tmp_ivl_38347 <= '0';
  tmp_ivl_38354 <= '0';
  tmp_ivl_38361 <= "00";
  tmp_ivl_38377 <= '0';
  tmp_ivl_38384 <= '0';
  tmp_ivl_38391 <= "00";
  tmp_ivl_3840 <= '0';
  tmp_ivl_38407 <= '0';
  tmp_ivl_38414 <= '0';
  tmp_ivl_38421 <= "00";
  tmp_ivl_38437 <= '0';
  tmp_ivl_38444 <= '0';
  tmp_ivl_38451 <= "00";
  tmp_ivl_38467 <= '0';
  tmp_ivl_38474 <= '0';
  tmp_ivl_38481 <= "00";
  tmp_ivl_38497 <= '0';
  tmp_ivl_38504 <= '0';
  tmp_ivl_38511 <= "00";
  tmp_ivl_38527 <= '0';
  tmp_ivl_38534 <= '0';
  tmp_ivl_38541 <= "00";
  tmp_ivl_38557 <= '0';
  tmp_ivl_3856 <= '0';
  tmp_ivl_38564 <= '0';
  tmp_ivl_38571 <= "00";
  tmp_ivl_38587 <= '0';
  tmp_ivl_38594 <= '0';
  tmp_ivl_386 <= '0';
  tmp_ivl_38601 <= "00";
  tmp_ivl_38617 <= '0';
  tmp_ivl_38624 <= '0';
  tmp_ivl_38631 <= "00";
  tmp_ivl_38647 <= '0';
  tmp_ivl_38654 <= '0';
  tmp_ivl_38661 <= "00";
  tmp_ivl_3867 <= '0';
  tmp_ivl_38677 <= '0';
  tmp_ivl_38684 <= '0';
  tmp_ivl_38691 <= "00";
  tmp_ivl_38707 <= '0';
  tmp_ivl_38714 <= '0';
  tmp_ivl_38721 <= "00";
  tmp_ivl_38737 <= '0';
  tmp_ivl_38744 <= '0';
  tmp_ivl_38751 <= "00";
  tmp_ivl_38767 <= '0';
  tmp_ivl_38774 <= '0';
  tmp_ivl_38781 <= "00";
  tmp_ivl_38797 <= '0';
  tmp_ivl_38804 <= '0';
  tmp_ivl_38811 <= "00";
  tmp_ivl_38827 <= '0';
  tmp_ivl_3883 <= '0';
  tmp_ivl_38834 <= '0';
  tmp_ivl_38841 <= "00";
  tmp_ivl_38857 <= '0';
  tmp_ivl_38864 <= '0';
  tmp_ivl_38871 <= "00";
  tmp_ivl_38887 <= '0';
  tmp_ivl_38894 <= '0';
  tmp_ivl_38901 <= "00";
  tmp_ivl_38917 <= '0';
  tmp_ivl_38924 <= '0';
  tmp_ivl_38931 <= "00";
  tmp_ivl_3894 <= '0';
  tmp_ivl_38947 <= '0';
  tmp_ivl_38954 <= '0';
  tmp_ivl_38961 <= "00";
  tmp_ivl_38977 <= '0';
  tmp_ivl_38984 <= '0';
  tmp_ivl_38991 <= "00";
  tmp_ivl_39007 <= '0';
  tmp_ivl_39014 <= '0';
  tmp_ivl_39021 <= "00";
  tmp_ivl_39037 <= '0';
  tmp_ivl_39044 <= '0';
  tmp_ivl_39051 <= "00";
  tmp_ivl_39067 <= '0';
  tmp_ivl_39074 <= '0';
  tmp_ivl_39081 <= "00";
  tmp_ivl_39097 <= '0';
  tmp_ivl_3910 <= '0';
  tmp_ivl_39104 <= '0';
  tmp_ivl_39111 <= "00";
  tmp_ivl_39127 <= '0';
  tmp_ivl_39134 <= '0';
  tmp_ivl_39141 <= "00";
  tmp_ivl_39157 <= '0';
  tmp_ivl_39164 <= '0';
  tmp_ivl_39171 <= "00";
  tmp_ivl_39187 <= '0';
  tmp_ivl_39194 <= '0';
  tmp_ivl_39201 <= "00";
  tmp_ivl_3921 <= '0';
  tmp_ivl_39217 <= '0';
  tmp_ivl_39224 <= '0';
  tmp_ivl_39231 <= "00";
  tmp_ivl_39247 <= '0';
  tmp_ivl_39254 <= '0';
  tmp_ivl_39261 <= "00";
  tmp_ivl_39277 <= '0';
  tmp_ivl_39284 <= '0';
  tmp_ivl_39291 <= "00";
  tmp_ivl_39307 <= '0';
  tmp_ivl_39314 <= '0';
  tmp_ivl_39321 <= "00";
  tmp_ivl_39337 <= '0';
  tmp_ivl_39344 <= '0';
  tmp_ivl_39351 <= "00";
  tmp_ivl_39367 <= '0';
  tmp_ivl_3937 <= '0';
  tmp_ivl_39374 <= '0';
  tmp_ivl_39381 <= "00";
  tmp_ivl_39397 <= '0';
  tmp_ivl_39404 <= '0';
  tmp_ivl_39411 <= "00";
  tmp_ivl_39427 <= '0';
  tmp_ivl_39434 <= '0';
  tmp_ivl_39441 <= "00";
  tmp_ivl_39457 <= '0';
  tmp_ivl_39464 <= '0';
  tmp_ivl_39471 <= "00";
  tmp_ivl_3948 <= '0';
  tmp_ivl_39487 <= '0';
  tmp_ivl_39494 <= '0';
  tmp_ivl_39501 <= "00";
  tmp_ivl_39517 <= '0';
  tmp_ivl_39524 <= '0';
  tmp_ivl_39531 <= "00";
  tmp_ivl_39547 <= '0';
  tmp_ivl_39554 <= '0';
  tmp_ivl_39561 <= "00";
  tmp_ivl_39577 <= '0';
  tmp_ivl_39584 <= '0';
  tmp_ivl_39591 <= "00";
  tmp_ivl_39607 <= '0';
  tmp_ivl_39614 <= '0';
  tmp_ivl_39621 <= "00";
  tmp_ivl_39637 <= '0';
  tmp_ivl_3964 <= '0';
  tmp_ivl_39644 <= '0';
  tmp_ivl_39651 <= "00";
  tmp_ivl_39667 <= '0';
  tmp_ivl_39674 <= '0';
  tmp_ivl_39681 <= "00";
  tmp_ivl_39697 <= '0';
  tmp_ivl_397 <= '0';
  tmp_ivl_39704 <= '0';
  tmp_ivl_39711 <= "00";
  tmp_ivl_39727 <= '0';
  tmp_ivl_39734 <= '0';
  tmp_ivl_39741 <= "00";
  tmp_ivl_3975 <= '0';
  tmp_ivl_39757 <= '0';
  tmp_ivl_39764 <= '0';
  tmp_ivl_39771 <= "00";
  tmp_ivl_39787 <= '0';
  tmp_ivl_39794 <= '0';
  tmp_ivl_39801 <= "00";
  tmp_ivl_39817 <= '0';
  tmp_ivl_39824 <= '0';
  tmp_ivl_39831 <= "00";
  tmp_ivl_39847 <= '0';
  tmp_ivl_39854 <= '0';
  tmp_ivl_39861 <= "00";
  tmp_ivl_39877 <= '0';
  tmp_ivl_39884 <= '0';
  tmp_ivl_39891 <= "00";
  tmp_ivl_39907 <= '0';
  tmp_ivl_3991 <= '0';
  tmp_ivl_39914 <= '0';
  tmp_ivl_39921 <= "00";
  tmp_ivl_39937 <= '0';
  tmp_ivl_39944 <= '0';
  tmp_ivl_39951 <= "00";
  tmp_ivl_39967 <= '0';
  tmp_ivl_39974 <= '0';
  tmp_ivl_39981 <= "00";
  tmp_ivl_39997 <= '0';
  tmp_ivl_40004 <= '0';
  tmp_ivl_40011 <= "00";
  tmp_ivl_4002 <= '0';
  tmp_ivl_40027 <= '0';
  tmp_ivl_40034 <= '0';
  tmp_ivl_40041 <= "00";
  tmp_ivl_40057 <= '0';
  tmp_ivl_40064 <= '0';
  tmp_ivl_40071 <= "00";
  tmp_ivl_40087 <= '0';
  tmp_ivl_40094 <= '0';
  tmp_ivl_40101 <= "00";
  tmp_ivl_40117 <= '0';
  tmp_ivl_40124 <= '0';
  tmp_ivl_40131 <= "00";
  tmp_ivl_40147 <= '0';
  tmp_ivl_40154 <= '0';
  tmp_ivl_40161 <= "00";
  tmp_ivl_40177 <= '0';
  tmp_ivl_4018 <= '0';
  tmp_ivl_40184 <= '0';
  tmp_ivl_40191 <= "00";
  tmp_ivl_40207 <= '0';
  tmp_ivl_40214 <= '0';
  tmp_ivl_40221 <= "00";
  tmp_ivl_40237 <= '0';
  tmp_ivl_40244 <= '0';
  tmp_ivl_40251 <= "00";
  tmp_ivl_40267 <= '0';
  tmp_ivl_40274 <= '0';
  tmp_ivl_40281 <= "00";
  tmp_ivl_4029 <= '0';
  tmp_ivl_40297 <= '0';
  tmp_ivl_40304 <= '0';
  tmp_ivl_40311 <= "00";
  tmp_ivl_40327 <= '0';
  tmp_ivl_40334 <= '0';
  tmp_ivl_40341 <= "00";
  tmp_ivl_40357 <= '0';
  tmp_ivl_40364 <= '0';
  tmp_ivl_40371 <= "00";
  tmp_ivl_40387 <= '0';
  tmp_ivl_40394 <= '0';
  tmp_ivl_40401 <= "00";
  tmp_ivl_40417 <= '0';
  tmp_ivl_40424 <= '0';
  tmp_ivl_40431 <= "00";
  tmp_ivl_40447 <= '0';
  tmp_ivl_4045 <= '0';
  tmp_ivl_40454 <= '0';
  tmp_ivl_40461 <= "00";
  tmp_ivl_40477 <= '0';
  tmp_ivl_40484 <= '0';
  tmp_ivl_40491 <= "00";
  tmp_ivl_40507 <= '0';
  tmp_ivl_40514 <= '0';
  tmp_ivl_40521 <= "00";
  tmp_ivl_40537 <= '0';
  tmp_ivl_40544 <= '0';
  tmp_ivl_40551 <= "00";
  tmp_ivl_4056 <= '0';
  tmp_ivl_40567 <= '0';
  tmp_ivl_40574 <= '0';
  tmp_ivl_40581 <= "00";
  tmp_ivl_40597 <= '0';
  tmp_ivl_40604 <= '0';
  tmp_ivl_40611 <= "00";
  tmp_ivl_40627 <= '0';
  tmp_ivl_40634 <= '0';
  tmp_ivl_40641 <= "00";
  tmp_ivl_40657 <= '0';
  tmp_ivl_40664 <= '0';
  tmp_ivl_40671 <= "00";
  tmp_ivl_40687 <= '0';
  tmp_ivl_40694 <= '0';
  tmp_ivl_40701 <= "00";
  tmp_ivl_40717 <= '0';
  tmp_ivl_4072 <= '0';
  tmp_ivl_40724 <= '0';
  tmp_ivl_40731 <= "00";
  tmp_ivl_40747 <= '0';
  tmp_ivl_40754 <= '0';
  tmp_ivl_40761 <= "00";
  tmp_ivl_40775 <= '0';
  tmp_ivl_40784 <= '0';
  tmp_ivl_40791 <= "00";
  tmp_ivl_40805 <= '0';
  tmp_ivl_40814 <= '0';
  tmp_ivl_40821 <= "00";
  tmp_ivl_4083 <= '0';
  tmp_ivl_40835 <= '0';
  tmp_ivl_40844 <= '0';
  tmp_ivl_40851 <= "00";
  tmp_ivl_40865 <= '0';
  tmp_ivl_40874 <= '0';
  tmp_ivl_40881 <= "00";
  tmp_ivl_40895 <= '0';
  tmp_ivl_40904 <= '0';
  tmp_ivl_40911 <= "00";
  tmp_ivl_40925 <= '0';
  tmp_ivl_40934 <= '0';
  tmp_ivl_40941 <= "00";
  tmp_ivl_40955 <= '0';
  tmp_ivl_40964 <= '0';
  tmp_ivl_40971 <= "00";
  tmp_ivl_40985 <= '0';
  tmp_ivl_4099 <= '0';
  tmp_ivl_40994 <= '0';
  tmp_ivl_41001 <= "00";
  tmp_ivl_41015 <= '0';
  tmp_ivl_41024 <= '0';
  tmp_ivl_41031 <= "00";
  tmp_ivl_41045 <= '0';
  tmp_ivl_41054 <= '0';
  tmp_ivl_41061 <= "00";
  tmp_ivl_41075 <= '0';
  tmp_ivl_41084 <= '0';
  tmp_ivl_41091 <= "00";
  tmp_ivl_4110 <= '0';
  tmp_ivl_41105 <= '0';
  tmp_ivl_41114 <= '0';
  tmp_ivl_41121 <= "00";
  tmp_ivl_41135 <= '0';
  tmp_ivl_41144 <= '0';
  tmp_ivl_41151 <= "00";
  tmp_ivl_41165 <= '0';
  tmp_ivl_41174 <= '0';
  tmp_ivl_41181 <= "00";
  tmp_ivl_41195 <= '0';
  tmp_ivl_41204 <= '0';
  tmp_ivl_41211 <= "00";
  tmp_ivl_41225 <= '0';
  tmp_ivl_41234 <= '0';
  tmp_ivl_41241 <= "00";
  tmp_ivl_41255 <= '0';
  tmp_ivl_4126 <= '0';
  tmp_ivl_41264 <= '0';
  tmp_ivl_41271 <= "00";
  tmp_ivl_41285 <= '0';
  tmp_ivl_41294 <= '0';
  tmp_ivl_41301 <= "00";
  tmp_ivl_41315 <= '0';
  tmp_ivl_41324 <= '0';
  tmp_ivl_41331 <= "00";
  tmp_ivl_41345 <= '0';
  tmp_ivl_41354 <= '0';
  tmp_ivl_41361 <= "00";
  tmp_ivl_4137 <= '0';
  tmp_ivl_41375 <= '0';
  tmp_ivl_41384 <= '0';
  tmp_ivl_41391 <= "00";
  tmp_ivl_41405 <= '0';
  tmp_ivl_41414 <= '0';
  tmp_ivl_41421 <= "00";
  tmp_ivl_41435 <= '0';
  tmp_ivl_41444 <= '0';
  tmp_ivl_41451 <= "00";
  tmp_ivl_41465 <= '0';
  tmp_ivl_41474 <= '0';
  tmp_ivl_41481 <= "00";
  tmp_ivl_41495 <= '0';
  tmp_ivl_415 <= '0';
  tmp_ivl_41504 <= '0';
  tmp_ivl_41511 <= "00";
  tmp_ivl_41525 <= '0';
  tmp_ivl_4153 <= '0';
  tmp_ivl_41534 <= '0';
  tmp_ivl_41541 <= "00";
  tmp_ivl_41555 <= '0';
  tmp_ivl_41564 <= '0';
  tmp_ivl_41571 <= "00";
  tmp_ivl_41585 <= '0';
  tmp_ivl_41594 <= '0';
  tmp_ivl_41601 <= "00";
  tmp_ivl_41615 <= '0';
  tmp_ivl_41624 <= '0';
  tmp_ivl_41631 <= "00";
  tmp_ivl_4164 <= '0';
  tmp_ivl_41645 <= '0';
  tmp_ivl_41654 <= '0';
  tmp_ivl_41661 <= "00";
  tmp_ivl_41675 <= '0';
  tmp_ivl_41684 <= '0';
  tmp_ivl_41691 <= "00";
  tmp_ivl_41705 <= '0';
  tmp_ivl_41714 <= '0';
  tmp_ivl_41721 <= "00";
  tmp_ivl_41735 <= '0';
  tmp_ivl_41744 <= '0';
  tmp_ivl_41751 <= "00";
  tmp_ivl_41765 <= '0';
  tmp_ivl_41774 <= '0';
  tmp_ivl_41781 <= "00";
  tmp_ivl_41795 <= '0';
  tmp_ivl_4180 <= '0';
  tmp_ivl_41804 <= '0';
  tmp_ivl_41811 <= "00";
  tmp_ivl_41825 <= '0';
  tmp_ivl_41834 <= '0';
  tmp_ivl_41841 <= "00";
  tmp_ivl_41855 <= '0';
  tmp_ivl_41864 <= '0';
  tmp_ivl_41871 <= "00";
  tmp_ivl_41885 <= '0';
  tmp_ivl_41894 <= '0';
  tmp_ivl_41901 <= "00";
  tmp_ivl_4191 <= '0';
  tmp_ivl_41915 <= '0';
  tmp_ivl_41922 <= '0';
  tmp_ivl_41929 <= "00";
  tmp_ivl_41943 <= '0';
  tmp_ivl_41950 <= '0';
  tmp_ivl_41957 <= "00";
  tmp_ivl_41971 <= '0';
  tmp_ivl_41978 <= '0';
  tmp_ivl_41985 <= "00";
  tmp_ivl_41999 <= '0';
  tmp_ivl_42006 <= '0';
  tmp_ivl_42013 <= "00";
  tmp_ivl_42027 <= '0';
  tmp_ivl_42034 <= '0';
  tmp_ivl_42041 <= "00";
  tmp_ivl_42055 <= '0';
  tmp_ivl_42062 <= '0';
  tmp_ivl_42069 <= "00";
  tmp_ivl_4207 <= '0';
  tmp_ivl_42083 <= '0';
  tmp_ivl_42090 <= '0';
  tmp_ivl_42097 <= "00";
  tmp_ivl_42111 <= '0';
  tmp_ivl_42118 <= '0';
  tmp_ivl_42125 <= "00";
  tmp_ivl_42139 <= '0';
  tmp_ivl_42146 <= '0';
  tmp_ivl_42153 <= "00";
  tmp_ivl_42167 <= '0';
  tmp_ivl_42174 <= '0';
  tmp_ivl_4218 <= '0';
  tmp_ivl_42181 <= "00";
  tmp_ivl_42197 <= '0';
  tmp_ivl_42204 <= '0';
  tmp_ivl_42211 <= "00";
  tmp_ivl_42225 <= '0';
  tmp_ivl_42232 <= '0';
  tmp_ivl_42239 <= "00";
  tmp_ivl_42255 <= '0';
  tmp_ivl_42262 <= '0';
  tmp_ivl_42269 <= "00";
  tmp_ivl_42283 <= '0';
  tmp_ivl_42290 <= '0';
  tmp_ivl_42297 <= "00";
  tmp_ivl_42311 <= '0';
  tmp_ivl_42318 <= '0';
  tmp_ivl_42325 <= "00";
  tmp_ivl_42339 <= '0';
  tmp_ivl_4234 <= '0';
  tmp_ivl_42346 <= '0';
  tmp_ivl_42353 <= "00";
  tmp_ivl_42367 <= '0';
  tmp_ivl_42374 <= '0';
  tmp_ivl_42381 <= "00";
  tmp_ivl_42395 <= '0';
  tmp_ivl_42402 <= '0';
  tmp_ivl_42409 <= "00";
  tmp_ivl_42423 <= '0';
  tmp_ivl_42430 <= '0';
  tmp_ivl_42437 <= "00";
  tmp_ivl_4245 <= '0';
  tmp_ivl_42451 <= '0';
  tmp_ivl_42458 <= '0';
  tmp_ivl_42465 <= "00";
  tmp_ivl_42479 <= '0';
  tmp_ivl_42486 <= '0';
  tmp_ivl_42493 <= "00";
  tmp_ivl_42507 <= '0';
  tmp_ivl_42514 <= '0';
  tmp_ivl_42521 <= "00";
  tmp_ivl_42535 <= '0';
  tmp_ivl_42542 <= '0';
  tmp_ivl_42549 <= "00";
  tmp_ivl_42563 <= '0';
  tmp_ivl_42570 <= '0';
  tmp_ivl_42577 <= "00";
  tmp_ivl_42591 <= '0';
  tmp_ivl_42598 <= '0';
  tmp_ivl_426 <= '0';
  tmp_ivl_42605 <= "00";
  tmp_ivl_4261 <= '0';
  tmp_ivl_42619 <= '0';
  tmp_ivl_42626 <= '0';
  tmp_ivl_42633 <= "00";
  tmp_ivl_42647 <= '0';
  tmp_ivl_42654 <= '0';
  tmp_ivl_42661 <= "00";
  tmp_ivl_42675 <= '0';
  tmp_ivl_42682 <= '0';
  tmp_ivl_42689 <= "00";
  tmp_ivl_42703 <= '0';
  tmp_ivl_42710 <= '0';
  tmp_ivl_42717 <= "00";
  tmp_ivl_4272 <= '0';
  tmp_ivl_42731 <= '0';
  tmp_ivl_42738 <= '0';
  tmp_ivl_42745 <= "00";
  tmp_ivl_42759 <= '0';
  tmp_ivl_42766 <= '0';
  tmp_ivl_42773 <= "00";
  tmp_ivl_42787 <= '0';
  tmp_ivl_42794 <= '0';
  tmp_ivl_42801 <= "00";
  tmp_ivl_42815 <= '0';
  tmp_ivl_42822 <= '0';
  tmp_ivl_42829 <= "00";
  tmp_ivl_42843 <= '0';
  tmp_ivl_42850 <= '0';
  tmp_ivl_42857 <= "00";
  tmp_ivl_42871 <= '0';
  tmp_ivl_42878 <= '0';
  tmp_ivl_4288 <= '0';
  tmp_ivl_42885 <= "00";
  tmp_ivl_42899 <= '0';
  tmp_ivl_42906 <= '0';
  tmp_ivl_42913 <= "00";
  tmp_ivl_42927 <= '0';
  tmp_ivl_42934 <= '0';
  tmp_ivl_42941 <= "00";
  tmp_ivl_42955 <= '0';
  tmp_ivl_42962 <= '0';
  tmp_ivl_42969 <= "00";
  tmp_ivl_42983 <= '0';
  tmp_ivl_4299 <= '0';
  tmp_ivl_42990 <= '0';
  tmp_ivl_42997 <= "00";
  tmp_ivl_43011 <= '0';
  tmp_ivl_43018 <= '0';
  tmp_ivl_43025 <= "00";
  tmp_ivl_43039 <= '0';
  tmp_ivl_43046 <= '0';
  tmp_ivl_43053 <= "00";
  tmp_ivl_43067 <= '0';
  tmp_ivl_43074 <= '0';
  tmp_ivl_43081 <= "00";
  tmp_ivl_43095 <= '0';
  tmp_ivl_43102 <= '0';
  tmp_ivl_43109 <= "00";
  tmp_ivl_43123 <= '0';
  tmp_ivl_43130 <= '0';
  tmp_ivl_43137 <= "00";
  tmp_ivl_4315 <= '0';
  tmp_ivl_43151 <= '0';
  tmp_ivl_43158 <= '0';
  tmp_ivl_43165 <= "00";
  tmp_ivl_43179 <= '0';
  tmp_ivl_43186 <= '0';
  tmp_ivl_43193 <= "00";
  tmp_ivl_43207 <= '0';
  tmp_ivl_43214 <= '0';
  tmp_ivl_43221 <= "00";
  tmp_ivl_43235 <= '0';
  tmp_ivl_43242 <= '0';
  tmp_ivl_43249 <= "00";
  tmp_ivl_4326 <= '0';
  tmp_ivl_43263 <= '0';
  tmp_ivl_43270 <= '0';
  tmp_ivl_43277 <= "00";
  tmp_ivl_43291 <= '0';
  tmp_ivl_43298 <= '0';
  tmp_ivl_43305 <= "00";
  tmp_ivl_43319 <= '0';
  tmp_ivl_43326 <= '0';
  tmp_ivl_43333 <= "00";
  tmp_ivl_43347 <= '0';
  tmp_ivl_43354 <= '0';
  tmp_ivl_43361 <= "00";
  tmp_ivl_43375 <= '0';
  tmp_ivl_43382 <= '0';
  tmp_ivl_43389 <= "00";
  tmp_ivl_43403 <= '0';
  tmp_ivl_43410 <= '0';
  tmp_ivl_43417 <= "00";
  tmp_ivl_4342 <= '0';
  tmp_ivl_43431 <= '0';
  tmp_ivl_43438 <= '0';
  tmp_ivl_43445 <= "00";
  tmp_ivl_43459 <= '0';
  tmp_ivl_43466 <= '0';
  tmp_ivl_43473 <= "00";
  tmp_ivl_43487 <= '0';
  tmp_ivl_43494 <= '0';
  tmp_ivl_43501 <= "00";
  tmp_ivl_43515 <= '0';
  tmp_ivl_43522 <= '0';
  tmp_ivl_43529 <= "00";
  tmp_ivl_4353 <= '0';
  tmp_ivl_43543 <= '0';
  tmp_ivl_43550 <= '0';
  tmp_ivl_43557 <= "00";
  tmp_ivl_43571 <= '0';
  tmp_ivl_43578 <= '0';
  tmp_ivl_43585 <= "00";
  tmp_ivl_43599 <= '0';
  tmp_ivl_43606 <= '0';
  tmp_ivl_43613 <= "00";
  tmp_ivl_43627 <= '0';
  tmp_ivl_43634 <= '0';
  tmp_ivl_43641 <= "00";
  tmp_ivl_43655 <= '0';
  tmp_ivl_43662 <= '0';
  tmp_ivl_43669 <= "00";
  tmp_ivl_43683 <= '0';
  tmp_ivl_4369 <= '0';
  tmp_ivl_43690 <= '0';
  tmp_ivl_43697 <= "00";
  tmp_ivl_43711 <= '0';
  tmp_ivl_43720 <= '0';
  tmp_ivl_43727 <= "00";
  tmp_ivl_43741 <= '0';
  tmp_ivl_43750 <= '0';
  tmp_ivl_43757 <= "00";
  tmp_ivl_43771 <= '0';
  tmp_ivl_43780 <= '0';
  tmp_ivl_43787 <= "00";
  tmp_ivl_4380 <= '0';
  tmp_ivl_43801 <= '0';
  tmp_ivl_43810 <= '0';
  tmp_ivl_43817 <= "00";
  tmp_ivl_43831 <= '0';
  tmp_ivl_43840 <= '0';
  tmp_ivl_43847 <= "00";
  tmp_ivl_43861 <= '0';
  tmp_ivl_43870 <= '0';
  tmp_ivl_43877 <= "00";
  tmp_ivl_43891 <= '0';
  tmp_ivl_43900 <= '0';
  tmp_ivl_43907 <= "00";
  tmp_ivl_43921 <= '0';
  tmp_ivl_43930 <= '0';
  tmp_ivl_43937 <= "00";
  tmp_ivl_43951 <= '0';
  tmp_ivl_4396 <= '0';
  tmp_ivl_43960 <= '0';
  tmp_ivl_43967 <= "00";
  tmp_ivl_43981 <= '0';
  tmp_ivl_43990 <= '0';
  tmp_ivl_43997 <= "00";
  tmp_ivl_44011 <= '0';
  tmp_ivl_44020 <= '0';
  tmp_ivl_44027 <= "00";
  tmp_ivl_44041 <= '0';
  tmp_ivl_44050 <= '0';
  tmp_ivl_44057 <= "00";
  tmp_ivl_4407 <= '0';
  tmp_ivl_44071 <= '0';
  tmp_ivl_44080 <= '0';
  tmp_ivl_44087 <= "00";
  tmp_ivl_44101 <= '0';
  tmp_ivl_44110 <= '0';
  tmp_ivl_44117 <= "00";
  tmp_ivl_44131 <= '0';
  tmp_ivl_44140 <= '0';
  tmp_ivl_44147 <= "00";
  tmp_ivl_44161 <= '0';
  tmp_ivl_44170 <= '0';
  tmp_ivl_44177 <= "00";
  tmp_ivl_44191 <= '0';
  tmp_ivl_44200 <= '0';
  tmp_ivl_44207 <= "00";
  tmp_ivl_44221 <= '0';
  tmp_ivl_4423 <= '0';
  tmp_ivl_44230 <= '0';
  tmp_ivl_44237 <= "00";
  tmp_ivl_44251 <= '0';
  tmp_ivl_44260 <= '0';
  tmp_ivl_44267 <= "00";
  tmp_ivl_44281 <= '0';
  tmp_ivl_44290 <= '0';
  tmp_ivl_44297 <= "00";
  tmp_ivl_44311 <= '0';
  tmp_ivl_44320 <= '0';
  tmp_ivl_44327 <= "00";
  tmp_ivl_4434 <= '0';
  tmp_ivl_44341 <= '0';
  tmp_ivl_44350 <= '0';
  tmp_ivl_44357 <= "00";
  tmp_ivl_44371 <= '0';
  tmp_ivl_44380 <= '0';
  tmp_ivl_44387 <= "00";
  tmp_ivl_444 <= '0';
  tmp_ivl_44401 <= '0';
  tmp_ivl_44410 <= '0';
  tmp_ivl_44417 <= "00";
  tmp_ivl_44431 <= '0';
  tmp_ivl_44440 <= '0';
  tmp_ivl_44447 <= "00";
  tmp_ivl_44461 <= '0';
  tmp_ivl_44470 <= '0';
  tmp_ivl_44477 <= "00";
  tmp_ivl_4450 <= '0';
  tmp_ivl_4461 <= '0';
  tmp_ivl_4477 <= '0';
  tmp_ivl_4488 <= '0';
  tmp_ivl_4504 <= '0';
  tmp_ivl_4515 <= '0';
  tmp_ivl_4531 <= '0';
  tmp_ivl_4542 <= '0';
  tmp_ivl_455 <= '0';
  tmp_ivl_4558 <= '0';
  tmp_ivl_4569 <= '0';
  tmp_ivl_4585 <= '0';
  tmp_ivl_4596 <= '0';
  tmp_ivl_4612 <= '0';
  tmp_ivl_4623 <= '0';
  tmp_ivl_4639 <= '0';
  tmp_ivl_4650 <= '0';
  tmp_ivl_4666 <= '0';
  tmp_ivl_4677 <= '0';
  tmp_ivl_4693 <= '0';
  tmp_ivl_4704 <= '0';
  tmp_ivl_4720 <= '0';
  tmp_ivl_473 <= '0';
  tmp_ivl_4731 <= '0';
  tmp_ivl_4747 <= '0';
  tmp_ivl_4758 <= '0';
  tmp_ivl_4774 <= '0';
  tmp_ivl_4785 <= '0';
  tmp_ivl_4801 <= '0';
  tmp_ivl_4812 <= '0';
  tmp_ivl_4828 <= '0';
  tmp_ivl_4839 <= '0';
  tmp_ivl_484 <= '0';
  tmp_ivl_4855 <= '0';
  tmp_ivl_4866 <= '0';
  tmp_ivl_4882 <= '0';
  tmp_ivl_4893 <= '0';
  tmp_ivl_49 <= '0';
  tmp_ivl_4909 <= '0';
  tmp_ivl_4920 <= '0';
  tmp_ivl_4936 <= '0';
  tmp_ivl_4947 <= '0';
  tmp_ivl_4963 <= '0';
  tmp_ivl_4974 <= '0';
  tmp_ivl_4990 <= '0';
  tmp_ivl_5001 <= '0';
  tmp_ivl_5017 <= '0';
  tmp_ivl_502 <= '0';
  tmp_ivl_5028 <= '0';
  tmp_ivl_5044 <= '0';
  tmp_ivl_5055 <= '0';
  tmp_ivl_5071 <= '0';
  tmp_ivl_5082 <= '0';
  tmp_ivl_5098 <= '0';
  tmp_ivl_5109 <= '0';
  tmp_ivl_5125 <= '0';
  tmp_ivl_513 <= '0';
  tmp_ivl_5136 <= '0';
  tmp_ivl_5152 <= '0';
  tmp_ivl_5163 <= '0';
  tmp_ivl_5179 <= '0';
  tmp_ivl_5190 <= '0';
  tmp_ivl_5206 <= '0';
  tmp_ivl_5217 <= '0';
  tmp_ivl_5233 <= '0';
  tmp_ivl_5244 <= '0';
  tmp_ivl_5260 <= '0';
  tmp_ivl_5271 <= '0';
  tmp_ivl_5287 <= '0';
  tmp_ivl_5298 <= '0';
  tmp_ivl_531 <= '0';
  tmp_ivl_5314 <= '0';
  tmp_ivl_5325 <= '0';
  tmp_ivl_5341 <= '0';
  tmp_ivl_5352 <= '0';
  tmp_ivl_5368 <= '0';
  tmp_ivl_5379 <= '0';
  tmp_ivl_5395 <= '0';
  tmp_ivl_5406 <= '0';
  tmp_ivl_542 <= '0';
  tmp_ivl_5422 <= '0';
  tmp_ivl_5433 <= '0';
  tmp_ivl_5449 <= '0';
  tmp_ivl_5460 <= '0';
  tmp_ivl_5476 <= '0';
  tmp_ivl_5487 <= '0';
  tmp_ivl_5503 <= '0';
  tmp_ivl_5514 <= '0';
  tmp_ivl_5530 <= '0';
  tmp_ivl_5541 <= '0';
  tmp_ivl_5557 <= '0';
  tmp_ivl_5568 <= '0';
  tmp_ivl_5584 <= '0';
  tmp_ivl_5595 <= '0';
  tmp_ivl_560 <= '0';
  tmp_ivl_5609 <= '0';
  tmp_ivl_5611 <= '0';
  tmp_ivl_5618 <= '0';
  tmp_ivl_5636 <= '0';
  tmp_ivl_5647 <= '0';
  tmp_ivl_5663 <= '0';
  tmp_ivl_5674 <= '0';
  tmp_ivl_5690 <= '0';
  tmp_ivl_5701 <= '0';
  tmp_ivl_571 <= '0';
  tmp_ivl_5717 <= '0';
  tmp_ivl_5728 <= '0';
  tmp_ivl_5735 <= '0';
  tmp_ivl_5744 <= '0';
  tmp_ivl_5751 <= '0';
  tmp_ivl_5767 <= '0';
  tmp_ivl_5778 <= '0';
  tmp_ivl_5798 <= '0';
  tmp_ivl_5809 <= '0';
  tmp_ivl_5816 <= '0';
  tmp_ivl_5823 <= '0';
  tmp_ivl_5830 <= '0';
  tmp_ivl_5848 <= '0';
  tmp_ivl_5859 <= '0';
  tmp_ivl_5873 <= '0';
  tmp_ivl_5875 <= '0';
  tmp_ivl_5882 <= '0';
  tmp_ivl_589 <= '0';
  tmp_ivl_5893 <= '0';
  tmp_ivl_5900 <= '0';
  tmp_ivl_5911 <= '0';
  tmp_ivl_5927 <= '0';
  tmp_ivl_5934 <= '0';
  tmp_ivl_5941 <= '0';
  tmp_ivl_5948 <= '0';
  tmp_ivl_5959 <= '0';
  tmp_ivl_5971 <= '0';
  tmp_ivl_5982 <= '0';
  tmp_ivl_5998 <= '0';
  tmp_ivl_600 <= '0';
  tmp_ivl_6009 <= '0';
  tmp_ivl_6016 <= '0';
  tmp_ivl_6023 <= '0';
  tmp_ivl_6030 <= '0';
  tmp_ivl_6046 <= '0';
  tmp_ivl_6057 <= '0';
  tmp_ivl_6064 <= '0';
  tmp_ivl_6071 <= '0';
  tmp_ivl_6078 <= '0';
  tmp_ivl_618 <= '0';
  tmp_ivl_629 <= '0';
  tmp_ivl_647 <= '0';
  tmp_ivl_658 <= '0';
  tmp_ivl_67 <= '0';
  tmp_ivl_676 <= '0';
  tmp_ivl_687 <= '0';
  tmp_ivl_705 <= '0';
  tmp_ivl_716 <= '0';
  tmp_ivl_734 <= '0';
  tmp_ivl_745 <= '0';
  tmp_ivl_763 <= '0';
  tmp_ivl_7694 <= '0';
  tmp_ivl_7703 <= '0';
  tmp_ivl_7719 <= '0';
  tmp_ivl_7726 <= '0';
  tmp_ivl_774 <= '0';
  tmp_ivl_7742 <= '0';
  tmp_ivl_7751 <= '0';
  tmp_ivl_7767 <= '0';
  tmp_ivl_7774 <= '0';
  tmp_ivl_7786 <= '0';
  tmp_ivl_7793 <= '0';
  tmp_ivl_78 <= '0';
  tmp_ivl_7809 <= '0';
  tmp_ivl_7818 <= '0';
  tmp_ivl_7834 <= '0';
  tmp_ivl_7841 <= '0';
  tmp_ivl_7853 <= '0';
  tmp_ivl_7860 <= '0';
  tmp_ivl_7880 <= '0';
  tmp_ivl_7889 <= '0';
  tmp_ivl_7905 <= '0';
  tmp_ivl_7912 <= '0';
  tmp_ivl_792 <= '0';
  tmp_ivl_7928 <= '0';
  tmp_ivl_7937 <= '0';
  tmp_ivl_7953 <= '0';
  tmp_ivl_7960 <= '0';
  tmp_ivl_7972 <= '0';
  tmp_ivl_7979 <= '0';
  tmp_ivl_7995 <= '0';
  tmp_ivl_8004 <= '0';
  tmp_ivl_8020 <= '0';
  tmp_ivl_8027 <= '0';
  tmp_ivl_803 <= '0';
  tmp_ivl_8039 <= '0';
  tmp_ivl_8046 <= '0';
  tmp_ivl_8066 <= '0';
  tmp_ivl_8075 <= '0';
  tmp_ivl_8091 <= '0';
  tmp_ivl_8098 <= '0';
  tmp_ivl_8114 <= '0';
  tmp_ivl_8123 <= '0';
  tmp_ivl_8139 <= '0';
  tmp_ivl_8146 <= '0';
  tmp_ivl_8158 <= '0';
  tmp_ivl_8165 <= '0';
  tmp_ivl_8181 <= '0';
  tmp_ivl_8190 <= '0';
  tmp_ivl_8206 <= '0';
  tmp_ivl_821 <= '0';
  tmp_ivl_8213 <= '0';
  tmp_ivl_8225 <= '0';
  tmp_ivl_8232 <= '0';
  tmp_ivl_8252 <= '0';
  tmp_ivl_8261 <= '0';
  tmp_ivl_8277 <= '0';
  tmp_ivl_8284 <= '0';
  tmp_ivl_8300 <= '0';
  tmp_ivl_8309 <= '0';
  tmp_ivl_832 <= '0';
  tmp_ivl_8325 <= '0';
  tmp_ivl_8332 <= '0';
  tmp_ivl_8344 <= '0';
  tmp_ivl_8351 <= '0';
  tmp_ivl_8367 <= '0';
  tmp_ivl_8376 <= '0';
  tmp_ivl_8392 <= '0';
  tmp_ivl_8399 <= '0';
  tmp_ivl_8411 <= '0';
  tmp_ivl_8418 <= '0';
  tmp_ivl_8438 <= '0';
  tmp_ivl_8447 <= '0';
  tmp_ivl_8463 <= '0';
  tmp_ivl_8470 <= '0';
  tmp_ivl_8486 <= '0';
  tmp_ivl_8495 <= '0';
  tmp_ivl_850 <= '0';
  tmp_ivl_8511 <= '0';
  tmp_ivl_8518 <= '0';
  tmp_ivl_8530 <= '0';
  tmp_ivl_8537 <= '0';
  tmp_ivl_8553 <= '0';
  tmp_ivl_8562 <= '0';
  tmp_ivl_8578 <= '0';
  tmp_ivl_8585 <= '0';
  tmp_ivl_8597 <= '0';
  tmp_ivl_8604 <= '0';
  tmp_ivl_861 <= '0';
  tmp_ivl_8624 <= '0';
  tmp_ivl_8633 <= '0';
  tmp_ivl_8649 <= '0';
  tmp_ivl_8656 <= '0';
  tmp_ivl_8672 <= '0';
  tmp_ivl_8681 <= '0';
  tmp_ivl_8697 <= '0';
  tmp_ivl_8704 <= '0';
  tmp_ivl_8716 <= '0';
  tmp_ivl_8723 <= '0';
  tmp_ivl_8739 <= '0';
  tmp_ivl_8748 <= '0';
  tmp_ivl_8764 <= '0';
  tmp_ivl_8771 <= '0';
  tmp_ivl_8783 <= '0';
  tmp_ivl_879 <= '0';
  tmp_ivl_8790 <= '0';
  tmp_ivl_8810 <= '0';
  tmp_ivl_8819 <= '0';
  tmp_ivl_8835 <= '0';
  tmp_ivl_8842 <= '0';
  tmp_ivl_8854 <= '0';
  tmp_ivl_8861 <= '0';
  tmp_ivl_8877 <= '0';
  tmp_ivl_8886 <= '0';
  tmp_ivl_890 <= '0';
  tmp_ivl_8902 <= '0';
  tmp_ivl_8909 <= '0';
  tmp_ivl_8921 <= '0';
  tmp_ivl_8928 <= '0';
  tmp_ivl_8948 <= '0';
  tmp_ivl_8957 <= '0';
  tmp_ivl_8973 <= '0';
  tmp_ivl_8980 <= '0';
  tmp_ivl_8996 <= '0';
  tmp_ivl_9 <= '0';
  tmp_ivl_9005 <= '0';
  tmp_ivl_9021 <= '0';
  tmp_ivl_9028 <= '0';
  tmp_ivl_9040 <= '0';
  tmp_ivl_9047 <= '0';
  tmp_ivl_9063 <= '0';
  tmp_ivl_9072 <= '0';
  tmp_ivl_908 <= '0';
  tmp_ivl_9088 <= '0';
  tmp_ivl_9095 <= '0';
  tmp_ivl_9107 <= '0';
  tmp_ivl_9114 <= '0';
  tmp_ivl_9134 <= '0';
  tmp_ivl_9143 <= '0';
  tmp_ivl_9159 <= '0';
  tmp_ivl_9166 <= '0';
  tmp_ivl_9178 <= '0';
  tmp_ivl_9185 <= '0';
  tmp_ivl_919 <= '0';
  tmp_ivl_9201 <= '0';
  tmp_ivl_9210 <= '0';
  tmp_ivl_9226 <= '0';
  tmp_ivl_9233 <= '0';
  tmp_ivl_9245 <= '0';
  tmp_ivl_9252 <= '0';
  tmp_ivl_9272 <= '0';
  tmp_ivl_9281 <= '0';
  tmp_ivl_9297 <= '0';
  tmp_ivl_9304 <= '0';
  tmp_ivl_9316 <= '0';
  tmp_ivl_9323 <= '0';
  tmp_ivl_9339 <= '0';
  tmp_ivl_9348 <= '0';
  tmp_ivl_9364 <= '0';
  tmp_ivl_937 <= '0';
  tmp_ivl_9371 <= '0';
  tmp_ivl_9383 <= '0';
  tmp_ivl_9390 <= '0';
  tmp_ivl_9410 <= '0';
  tmp_ivl_9419 <= '0';
  tmp_ivl_9435 <= '0';
  tmp_ivl_9442 <= '0';
  tmp_ivl_9454 <= '0';
  tmp_ivl_9461 <= '0';
  tmp_ivl_9477 <= '0';
  tmp_ivl_948 <= '0';
  tmp_ivl_9486 <= '0';
  tmp_ivl_9502 <= '0';
  tmp_ivl_9509 <= '0';
  tmp_ivl_9521 <= '0';
  tmp_ivl_9528 <= '0';
  tmp_ivl_9548 <= '0';
  tmp_ivl_9557 <= '0';
  tmp_ivl_9573 <= '0';
  tmp_ivl_9580 <= '0';
  tmp_ivl_9592 <= '0';
  tmp_ivl_9599 <= '0';
  tmp_ivl_96 <= '0';
  tmp_ivl_9615 <= '0';
  tmp_ivl_9624 <= '0';
  tmp_ivl_9640 <= '0';
  tmp_ivl_9647 <= '0';
  tmp_ivl_9659 <= '0';
  tmp_ivl_966 <= '0';
  tmp_ivl_9666 <= '0';
  tmp_ivl_9682 <= '0';
  tmp_ivl_9689 <= '0';
  tmp_ivl_9705 <= '0';
  tmp_ivl_9714 <= '0';
  tmp_ivl_9730 <= '0';
  tmp_ivl_9737 <= '0';
  tmp_ivl_9749 <= '0';
  tmp_ivl_9756 <= '0';
  tmp_ivl_977 <= '0';
  tmp_ivl_9772 <= '0';
  tmp_ivl_9779 <= '0';
  tmp_ivl_9795 <= '0';
  tmp_ivl_9804 <= '0';
  tmp_ivl_9820 <= '0';
  tmp_ivl_9827 <= '0';
  tmp_ivl_9839 <= '0';
  tmp_ivl_9846 <= '0';
  tmp_ivl_9866 <= '0';
  tmp_ivl_9875 <= '0';
  tmp_ivl_9891 <= '0';
  tmp_ivl_9898 <= '0';
  tmp_ivl_9910 <= '0';
  tmp_ivl_9917 <= '0';
  tmp_ivl_9933 <= '0';
  tmp_ivl_9942 <= '0';
  tmp_ivl_995 <= '0';
  tmp_ivl_9958 <= '0';
  tmp_ivl_9965 <= '0';
  tmp_ivl_9977 <= '0';
  tmp_ivl_9984 <= '0';
end architecture;
